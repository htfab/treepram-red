magic
tech sky130A
magscale 1 2
timestamp 1636885634
<< locali >>
rect 97917 637687 97951 637925
rect 117145 637823 117179 637925
rect 473369 637755 473403 638265
rect 502533 637619 502567 638265
rect 523325 636871 523359 638265
rect 75101 62135 75135 63189
rect 78505 62883 78539 62985
rect 497565 62815 497599 63189
rect 108313 3927 108347 4097
rect 69673 3791 69707 3893
rect 98653 3791 98687 3893
rect 65349 3757 65533 3791
rect 34621 3383 34655 3621
rect 52469 2975 52503 3689
rect 65349 3655 65383 3757
rect 69305 3655 69339 3757
rect 57161 3315 57195 3485
rect 61577 2839 61611 3145
rect 79333 2975 79367 3757
rect 344661 3587 344695 3825
rect 84393 2975 84427 3213
rect 91109 2907 91143 3349
rect 93869 3247 93903 3417
rect 439421 3383 439455 3961
rect 451105 3043 451139 4097
rect 452485 3791 452519 4029
rect 452577 3791 452611 3893
rect 456625 3859 456659 4029
rect 462087 3689 462329 3723
rect 465917 3587 465951 3757
rect 502901 3315 502935 3621
rect 514033 3179 514067 3281
rect 535009 3179 535043 3553
rect 468769 2907 468803 3077
rect 542277 3043 542311 3145
rect 542277 3009 542553 3043
rect 518449 2907 518483 3009
rect 542921 2907 542955 3281
rect 546877 2975 546911 3349
rect 582389 3043 582423 62781
<< viali >>
rect 473369 638265 473403 638299
rect 97917 637925 97951 637959
rect 117145 637925 117179 637959
rect 117145 637789 117179 637823
rect 473369 637721 473403 637755
rect 502533 638265 502567 638299
rect 97917 637653 97951 637687
rect 502533 637585 502567 637619
rect 523325 638265 523359 638299
rect 523325 636837 523359 636871
rect 75101 63189 75135 63223
rect 497565 63189 497599 63223
rect 78505 62985 78539 63019
rect 78505 62849 78539 62883
rect 497565 62781 497599 62815
rect 582389 62781 582423 62815
rect 75101 62101 75135 62135
rect 108313 4097 108347 4131
rect 451105 4097 451139 4131
rect 69673 3893 69707 3927
rect 98653 3893 98687 3927
rect 108313 3893 108347 3927
rect 439421 3961 439455 3995
rect 65533 3757 65567 3791
rect 69305 3757 69339 3791
rect 69673 3757 69707 3791
rect 79333 3757 79367 3791
rect 98653 3757 98687 3791
rect 344661 3825 344695 3859
rect 52469 3689 52503 3723
rect 34621 3621 34655 3655
rect 34621 3349 34655 3383
rect 65349 3621 65383 3655
rect 69305 3621 69339 3655
rect 57161 3485 57195 3519
rect 57161 3281 57195 3315
rect 52469 2941 52503 2975
rect 61577 3145 61611 3179
rect 344661 3553 344695 3587
rect 93869 3417 93903 3451
rect 91109 3349 91143 3383
rect 79333 2941 79367 2975
rect 84393 3213 84427 3247
rect 84393 2941 84427 2975
rect 439421 3349 439455 3383
rect 93869 3213 93903 3247
rect 452485 4029 452519 4063
rect 456625 4029 456659 4063
rect 452485 3757 452519 3791
rect 452577 3893 452611 3927
rect 456625 3825 456659 3859
rect 452577 3757 452611 3791
rect 465917 3757 465951 3791
rect 462053 3689 462087 3723
rect 462329 3689 462363 3723
rect 465917 3553 465951 3587
rect 502901 3621 502935 3655
rect 535009 3553 535043 3587
rect 502901 3281 502935 3315
rect 514033 3281 514067 3315
rect 514033 3145 514067 3179
rect 546877 3349 546911 3383
rect 542921 3281 542955 3315
rect 535009 3145 535043 3179
rect 542277 3145 542311 3179
rect 451105 3009 451139 3043
rect 468769 3077 468803 3111
rect 91109 2873 91143 2907
rect 468769 2873 468803 2907
rect 518449 3009 518483 3043
rect 542553 3009 542587 3043
rect 518449 2873 518483 2907
rect 582389 3009 582423 3043
rect 546877 2941 546911 2975
rect 542921 2873 542955 2907
rect 61577 2805 61611 2839
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 327074 700992 327080 701004
rect 154172 700964 327080 700992
rect 154172 700952 154178 700964
rect 327074 700952 327080 700964
rect 327132 700952 327138 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 322934 700924 322940 700936
rect 137888 700896 322940 700924
rect 137888 700884 137894 700896
rect 322934 700884 322940 700896
rect 322992 700884 322998 700936
rect 260742 700816 260748 700868
rect 260800 700856 260806 700868
rect 462314 700856 462320 700868
rect 260800 700828 462320 700856
rect 260800 700816 260806 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 264882 700748 264888 700800
rect 264940 700788 264946 700800
rect 478506 700788 478512 700800
rect 264940 700760 478512 700788
rect 264940 700748 264946 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 339494 700720 339500 700732
rect 89220 700692 339500 700720
rect 89220 700680 89226 700692
rect 339494 700680 339500 700692
rect 339552 700680 339558 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 335354 700652 335360 700664
rect 73028 700624 335360 700652
rect 73028 700612 73034 700624
rect 335354 700612 335360 700624
rect 335412 700612 335418 700664
rect 342898 700612 342904 700664
rect 342956 700652 342962 700664
rect 364978 700652 364984 700664
rect 342956 700624 364984 700652
rect 342956 700612 342962 700624
rect 364978 700612 364984 700624
rect 365036 700612 365042 700664
rect 248322 700544 248328 700596
rect 248380 700584 248386 700596
rect 527174 700584 527180 700596
rect 248380 700556 527180 700584
rect 248380 700544 248386 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 166258 700516 166264 700528
rect 105504 700488 166264 700516
rect 105504 700476 105510 700488
rect 166258 700476 166264 700488
rect 166316 700476 166322 700528
rect 235166 700476 235172 700528
rect 235224 700516 235230 700528
rect 242158 700516 242164 700528
rect 235224 700488 242164 700516
rect 235224 700476 235230 700488
rect 242158 700476 242164 700488
rect 242216 700476 242222 700528
rect 252462 700476 252468 700528
rect 252520 700516 252526 700528
rect 543458 700516 543464 700528
rect 252520 700488 543464 700516
rect 252520 700476 252526 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 343634 700448 343640 700460
rect 40552 700420 343640 700448
rect 40552 700408 40558 700420
rect 343634 700408 343640 700420
rect 343692 700408 343698 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 351914 700380 351920 700392
rect 24360 700352 351920 700380
rect 24360 700340 24366 700352
rect 351914 700340 351920 700352
rect 351972 700340 351978 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 347866 700312 347872 700324
rect 8168 700284 347872 700312
rect 8168 700272 8174 700284
rect 347866 700272 347872 700284
rect 347924 700272 347930 700324
rect 349798 700272 349804 700324
rect 349856 700312 349862 700324
rect 429838 700312 429844 700324
rect 349856 700284 429844 700312
rect 349856 700272 349862 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 457438 700272 457444 700324
rect 457496 700312 457502 700324
rect 494790 700312 494796 700324
rect 457496 700284 494796 700312
rect 457496 700272 457502 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 526438 700272 526444 700324
rect 526496 700312 526502 700324
rect 559650 700312 559656 700324
rect 526496 700284 559656 700312
rect 526496 700272 526502 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 277302 700204 277308 700256
rect 277360 700244 277366 700256
rect 413646 700244 413652 700256
rect 277360 700216 413652 700244
rect 277360 700204 277366 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 273162 700136 273168 700188
rect 273220 700176 273226 700188
rect 397454 700176 397460 700188
rect 273220 700148 397460 700176
rect 273220 700136 273226 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 310514 700108 310520 700120
rect 202840 700080 310520 700108
rect 202840 700068 202846 700080
rect 310514 700068 310520 700080
rect 310572 700068 310578 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 314654 700040 314660 700052
rect 219032 700012 314660 700040
rect 219032 700000 219038 700012
rect 314654 700000 314660 700012
rect 314712 700000 314718 700052
rect 289722 699932 289728 699984
rect 289780 699972 289786 699984
rect 348786 699972 348792 699984
rect 289780 699944 348792 699972
rect 289780 699932 289786 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 285582 699864 285588 699916
rect 285640 699904 285646 699916
rect 332502 699904 332508 699916
rect 285640 699876 332508 699904
rect 285640 699864 285646 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 298094 699836 298100 699848
rect 267700 699808 298100 699836
rect 267700 699796 267706 699808
rect 298094 699796 298100 699808
rect 298152 699796 298158 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 302234 699768 302240 699780
rect 283892 699740 302240 699768
rect 283892 699728 283898 699740
rect 302234 699728 302240 699740
rect 302292 699728 302298 699780
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235902 696940 235908 696992
rect 235960 696980 235966 696992
rect 580166 696980 580172 696992
rect 235960 696952 580172 696980
rect 235960 696940 235966 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 240042 683204 240048 683256
rect 240100 683244 240106 683256
rect 580166 683244 580172 683256
rect 240100 683216 580172 683244
rect 240100 683204 240106 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 356054 683176 356060 683188
rect 3476 683148 356060 683176
rect 3476 683136 3482 683148
rect 356054 683136 356060 683148
rect 356112 683136 356118 683188
rect 231762 670760 231768 670812
rect 231820 670800 231826 670812
rect 580166 670800 580172 670812
rect 231820 670772 580172 670800
rect 231820 670760 231826 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 364334 670732 364340 670744
rect 3568 670704 364340 670732
rect 3568 670692 3574 670704
rect 364334 670692 364340 670704
rect 364392 670692 364398 670744
rect 242158 668584 242164 668636
rect 242216 668624 242222 668636
rect 306374 668624 306380 668636
rect 242216 668596 306380 668624
rect 242216 668584 242222 668596
rect 306374 668584 306380 668596
rect 306432 668584 306438 668636
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 360194 656928 360200 656940
rect 3476 656900 360200 656928
rect 3476 656888 3482 656900
rect 360194 656888 360200 656900
rect 360252 656888 360258 656940
rect 256326 643696 256332 643748
rect 256384 643736 256390 643748
rect 457438 643736 457444 643748
rect 256384 643708 457444 643736
rect 256384 643696 256390 643708
rect 457438 643696 457444 643708
rect 457496 643696 457502 643748
rect 222930 643084 222936 643136
rect 222988 643124 222994 643136
rect 580166 643124 580172 643136
rect 222988 643096 580172 643124
rect 222988 643084 222994 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 293954 642676 293960 642728
rect 294012 642716 294018 642728
rect 299474 642716 299480 642728
rect 294012 642688 299480 642716
rect 294012 642676 294018 642688
rect 299474 642676 299480 642688
rect 299532 642676 299538 642728
rect 281350 642608 281356 642660
rect 281408 642648 281414 642660
rect 342898 642648 342904 642660
rect 281408 642620 342904 642648
rect 281408 642608 281414 642620
rect 342898 642608 342904 642620
rect 342956 642608 342962 642660
rect 268838 642540 268844 642592
rect 268896 642580 268902 642592
rect 349798 642580 349804 642592
rect 268896 642552 349804 642580
rect 268896 642540 268902 642552
rect 349798 642540 349804 642552
rect 349856 642540 349862 642592
rect 171042 642472 171048 642524
rect 171100 642512 171106 642524
rect 318978 642512 318984 642524
rect 171100 642484 318984 642512
rect 171100 642472 171106 642484
rect 318978 642472 318984 642484
rect 319036 642472 319042 642524
rect 166258 642404 166264 642456
rect 166316 642444 166322 642456
rect 331490 642444 331496 642456
rect 166316 642416 331496 642444
rect 166316 642404 166322 642416
rect 331490 642404 331496 642416
rect 331548 642404 331554 642456
rect 243814 642336 243820 642388
rect 243872 642376 243878 642388
rect 526438 642376 526444 642388
rect 243872 642348 526444 642376
rect 243872 642336 243878 642348
rect 526438 642336 526444 642348
rect 526496 642336 526502 642388
rect 32398 641656 32404 641708
rect 32456 641696 32462 641708
rect 486050 641696 486056 641708
rect 32456 641668 486056 641696
rect 32456 641656 32462 641668
rect 486050 641656 486056 641668
rect 486108 641656 486114 641708
rect 176930 641588 176936 641640
rect 176988 641628 176994 641640
rect 369854 641628 369860 641640
rect 176988 641600 369860 641628
rect 176988 641588 176994 641600
rect 369854 641588 369860 641600
rect 369912 641588 369918 641640
rect 43530 641520 43536 641572
rect 43588 641560 43594 641572
rect 390002 641560 390008 641572
rect 43588 641532 390008 641560
rect 43588 641520 43594 641532
rect 390002 641520 390008 641532
rect 390060 641520 390066 641572
rect 189442 641452 189448 641504
rect 189500 641492 189506 641504
rect 536098 641492 536104 641504
rect 189500 641464 536104 641492
rect 189500 641452 189506 641464
rect 536098 641452 536104 641464
rect 536156 641452 536162 641504
rect 214558 641384 214564 641436
rect 214616 641424 214622 641436
rect 569310 641424 569316 641436
rect 214616 641396 569316 641424
rect 214616 641384 214622 641396
rect 569310 641384 569316 641396
rect 569368 641384 569374 641436
rect 139394 641316 139400 641368
rect 139452 641356 139458 641368
rect 189074 641356 189080 641368
rect 139452 641328 189080 641356
rect 139452 641316 139458 641328
rect 189074 641316 189080 641328
rect 189132 641316 189138 641368
rect 202046 641316 202052 641368
rect 202104 641356 202110 641368
rect 558270 641356 558276 641368
rect 202104 641328 558276 641356
rect 202104 641316 202110 641328
rect 558270 641316 558276 641328
rect 558328 641316 558334 641368
rect 50430 641248 50436 641300
rect 50488 641288 50494 641300
rect 423398 641288 423404 641300
rect 50488 641260 423404 641288
rect 50488 641248 50494 641260
rect 423398 641248 423404 641260
rect 423456 641248 423462 641300
rect 53190 641180 53196 641232
rect 53248 641220 53254 641232
rect 435910 641220 435916 641232
rect 53248 641192 435916 641220
rect 53248 641180 53254 641192
rect 435910 641180 435916 641192
rect 435968 641180 435974 641232
rect 168558 641112 168564 641164
rect 168616 641152 168622 641164
rect 551370 641152 551376 641164
rect 168616 641124 551376 641152
rect 168616 641112 168622 641124
rect 551370 641112 551376 641124
rect 551428 641112 551434 641164
rect 14458 641044 14464 641096
rect 14516 641084 14522 641096
rect 402514 641084 402520 641096
rect 14516 641056 402520 641084
rect 14516 641044 14522 641056
rect 402514 641044 402520 641056
rect 402572 641044 402578 641096
rect 415854 641044 415860 641096
rect 415912 641084 415918 641096
rect 477678 641084 477684 641096
rect 415912 641056 477684 641084
rect 415912 641044 415918 641056
rect 477678 641044 477684 641056
rect 477736 641044 477742 641096
rect 172790 640976 172796 641028
rect 172848 641016 172854 641028
rect 562318 641016 562324 641028
rect 172848 640988 562324 641016
rect 172848 640976 172854 640988
rect 562318 640976 562324 640988
rect 562376 640976 562382 641028
rect 40678 640908 40684 640960
rect 40736 640948 40742 640960
rect 440142 640948 440148 640960
rect 40736 640920 440148 640948
rect 40736 640908 40742 640920
rect 440142 640908 440148 640920
rect 440200 640908 440206 640960
rect 15838 640840 15844 640892
rect 15896 640880 15902 640892
rect 415026 640880 415032 640892
rect 15896 640852 415032 640880
rect 15896 640840 15902 640852
rect 415026 640840 415032 640852
rect 415084 640840 415090 640892
rect 435358 640840 435364 640892
rect 435416 640880 435422 640892
rect 527818 640880 527824 640892
rect 435416 640852 527824 640880
rect 435416 640840 435422 640852
rect 527818 640840 527824 640852
rect 527876 640840 527882 640892
rect 50338 640772 50344 640824
rect 50396 640812 50402 640824
rect 452654 640812 452660 640824
rect 50396 640784 452660 640812
rect 50396 640772 50402 640784
rect 452654 640772 452660 640784
rect 452712 640772 452718 640824
rect 143534 640704 143540 640756
rect 143592 640744 143598 640756
rect 547230 640744 547236 640756
rect 143592 640716 547236 640744
rect 143592 640704 143598 640716
rect 547230 640704 547236 640716
rect 547288 640704 547294 640756
rect 51718 640636 51724 640688
rect 51776 640676 51782 640688
rect 461026 640676 461032 640688
rect 51776 640648 461032 640676
rect 51776 640636 51782 640648
rect 461026 640636 461032 640648
rect 461084 640636 461090 640688
rect 118510 640568 118516 640620
rect 118568 640608 118574 640620
rect 542998 640608 543004 640620
rect 118568 640580 543004 640608
rect 118568 640568 118574 640580
rect 542998 640568 543004 640580
rect 543056 640568 543062 640620
rect 105906 640500 105912 640552
rect 105964 640540 105970 640552
rect 531958 640540 531964 640552
rect 105964 640512 531964 640540
rect 105964 640500 105970 640512
rect 531958 640500 531964 640512
rect 532016 640500 532022 640552
rect 53098 640432 53104 640484
rect 53156 640472 53162 640484
rect 490190 640472 490196 640484
rect 53156 640444 490196 640472
rect 53156 640432 53162 640444
rect 490190 640432 490196 640444
rect 490248 640432 490254 640484
rect 18598 640364 18604 640416
rect 18656 640404 18662 640416
rect 465166 640404 465172 640416
rect 18656 640376 465172 640404
rect 18656 640364 18662 640376
rect 465166 640364 465172 640376
rect 465224 640364 465230 640416
rect 164418 640296 164424 640348
rect 164476 640336 164482 640348
rect 175918 640336 175924 640348
rect 164476 640308 175924 640336
rect 164476 640296 164482 640308
rect 175918 640296 175924 640308
rect 175976 640296 175982 640348
rect 218698 640228 218704 640280
rect 218756 640268 218762 640280
rect 538950 640268 538956 640280
rect 218756 640240 538956 640268
rect 218756 640228 218762 640240
rect 538950 640228 538956 640240
rect 539008 640228 539014 640280
rect 206186 640160 206192 640212
rect 206244 640200 206250 640212
rect 537570 640200 537576 640212
rect 206244 640172 537576 640200
rect 206244 640160 206250 640172
rect 537570 640160 537576 640172
rect 537628 640160 537634 640212
rect 193674 640092 193680 640144
rect 193732 640132 193738 640144
rect 536190 640132 536196 640144
rect 193732 640104 536196 640132
rect 193732 640092 193738 640104
rect 536190 640092 536196 640104
rect 536248 640092 536254 640144
rect 181162 640024 181168 640076
rect 181220 640064 181226 640076
rect 533430 640064 533436 640076
rect 181220 640036 533436 640064
rect 181220 640024 181226 640036
rect 533430 640024 533436 640036
rect 533488 640024 533494 640076
rect 7650 639956 7656 640008
rect 7708 639996 7714 640008
rect 369118 639996 369124 640008
rect 7708 639968 369124 639996
rect 7708 639956 7714 639968
rect 369118 639956 369124 639968
rect 369176 639956 369182 640008
rect 369854 639956 369860 640008
rect 369912 639996 369918 640008
rect 580442 639996 580448 640008
rect 369912 639968 580448 639996
rect 369912 639956 369918 639968
rect 580442 639956 580448 639968
rect 580500 639956 580506 640008
rect 11790 639888 11796 639940
rect 11848 639928 11854 639940
rect 381630 639928 381636 639940
rect 11848 639900 381636 639928
rect 11848 639888 11854 639900
rect 381630 639888 381636 639900
rect 381688 639888 381694 639940
rect 14550 639820 14556 639872
rect 14608 639860 14614 639872
rect 394142 639860 394148 639872
rect 14608 639832 394148 639860
rect 14608 639820 14614 639832
rect 394142 639820 394148 639832
rect 394200 639820 394206 639872
rect 15930 639752 15936 639804
rect 15988 639792 15994 639804
rect 406654 639792 406660 639804
rect 15988 639764 406660 639792
rect 15988 639752 15994 639764
rect 406654 639752 406660 639764
rect 406712 639752 406718 639804
rect 156046 639684 156052 639736
rect 156104 639724 156110 639736
rect 548610 639724 548616 639736
rect 156104 639696 548616 639724
rect 156104 639684 156110 639696
rect 548610 639684 548616 639696
rect 548668 639684 548674 639736
rect 17310 639616 17316 639668
rect 17368 639656 17374 639668
rect 419258 639656 419264 639668
rect 17368 639628 419264 639656
rect 17368 639616 17374 639628
rect 419258 639616 419264 639628
rect 419316 639616 419322 639668
rect 18690 639548 18696 639600
rect 18748 639588 18754 639600
rect 431770 639588 431776 639600
rect 18748 639560 431776 639588
rect 18748 639548 18754 639560
rect 431770 639548 431776 639560
rect 431828 639548 431834 639600
rect 131022 639480 131028 639532
rect 131080 639520 131086 639532
rect 544470 639520 544476 639532
rect 131080 639492 544476 639520
rect 131080 639480 131086 639492
rect 544470 639480 544476 639492
rect 544528 639480 544534 639532
rect 21450 639412 21456 639464
rect 21508 639452 21514 639464
rect 444282 639452 444288 639464
rect 21508 639424 444288 639452
rect 21508 639412 21514 639424
rect 444282 639412 444288 639424
rect 444340 639412 444346 639464
rect 22738 639344 22744 639396
rect 22796 639384 22802 639396
rect 456794 639384 456800 639396
rect 22796 639356 456800 639384
rect 22796 639344 22802 639356
rect 456794 639344 456800 639356
rect 456852 639344 456858 639396
rect 93394 639276 93400 639328
rect 93452 639316 93458 639328
rect 530578 639316 530584 639328
rect 93452 639288 530584 639316
rect 93452 639276 93458 639288
rect 530578 639276 530584 639288
rect 530636 639276 530642 639328
rect 25498 639208 25504 639260
rect 25556 639248 25562 639260
rect 469306 639248 469312 639260
rect 25556 639220 469312 639248
rect 25556 639208 25562 639220
rect 469306 639208 469312 639220
rect 469364 639208 469370 639260
rect 36538 639140 36544 639192
rect 36596 639180 36602 639192
rect 481910 639180 481916 639192
rect 36596 639152 481916 639180
rect 36596 639140 36602 639152
rect 481910 639140 481916 639152
rect 481968 639140 481974 639192
rect 39298 639072 39304 639124
rect 39356 639112 39362 639124
rect 494422 639112 494428 639124
rect 39356 639084 494428 639112
rect 39356 639072 39362 639084
rect 494422 639072 494428 639084
rect 494480 639072 494486 639124
rect 47578 639004 47584 639056
rect 47636 639044 47642 639056
rect 506934 639044 506940 639056
rect 47636 639016 506940 639044
rect 47636 639004 47642 639016
rect 506934 639004 506940 639016
rect 506992 639004 506998 639056
rect 80882 638936 80888 638988
rect 80940 638976 80946 638988
rect 540238 638976 540244 638988
rect 80940 638948 540244 638976
rect 80940 638936 80946 638948
rect 540238 638936 540244 638948
rect 540296 638936 540302 638988
rect 227070 638868 227076 638920
rect 227128 638908 227134 638920
rect 530670 638908 530676 638920
rect 227128 638880 530676 638908
rect 227128 638868 227134 638880
rect 530670 638868 530676 638880
rect 530728 638868 530734 638920
rect 189074 638800 189080 638852
rect 189132 638840 189138 638852
rect 580258 638840 580264 638852
rect 189132 638812 580264 638840
rect 189132 638800 189138 638812
rect 580258 638800 580264 638812
rect 580316 638800 580322 638852
rect 40862 638732 40868 638784
rect 40920 638772 40926 638784
rect 377490 638772 377496 638784
rect 40920 638744 377496 638772
rect 40920 638732 40926 638744
rect 377490 638732 377496 638744
rect 377548 638732 377554 638784
rect 175918 638664 175924 638716
rect 175976 638704 175982 638716
rect 580350 638704 580356 638716
rect 175976 638676 580356 638704
rect 175976 638664 175982 638676
rect 580350 638664 580356 638676
rect 580408 638664 580414 638716
rect 3510 638596 3516 638648
rect 3568 638636 3574 638648
rect 415854 638636 415860 638648
rect 3568 638608 415860 638636
rect 3568 638596 3574 638608
rect 415854 638596 415860 638608
rect 415912 638596 415918 638648
rect 160554 638528 160560 638580
rect 160612 638568 160618 638580
rect 537478 638568 537484 638580
rect 160612 638540 537484 638568
rect 160612 638528 160618 638540
rect 537478 638528 537484 638540
rect 537536 638528 537542 638580
rect 152274 638460 152280 638512
rect 152332 638500 152338 638512
rect 532050 638500 532056 638512
rect 152332 638472 532056 638500
rect 152332 638460 152338 638472
rect 532050 638460 532056 638472
rect 532108 638460 532114 638512
rect 43438 638392 43444 638444
rect 43496 638432 43502 638444
rect 448054 638432 448060 638444
rect 43496 638404 448060 638432
rect 43496 638392 43502 638404
rect 448054 638392 448060 638404
rect 448112 638392 448118 638444
rect 135254 638324 135260 638376
rect 135312 638364 135318 638376
rect 538858 638364 538864 638376
rect 135312 638336 538864 638364
rect 135312 638324 135318 638336
rect 538858 638324 538864 638336
rect 538916 638324 538922 638376
rect 17218 638256 17224 638308
rect 17276 638296 17282 638308
rect 427262 638296 427268 638308
rect 17276 638268 427268 638296
rect 17276 638256 17282 638268
rect 427262 638256 427268 638268
rect 427320 638256 427326 638308
rect 473354 638296 473360 638308
rect 473315 638268 473360 638296
rect 473354 638256 473360 638268
rect 473412 638256 473418 638308
rect 502518 638296 502524 638308
rect 502479 638268 502524 638296
rect 502518 638256 502524 638268
rect 502576 638256 502582 638308
rect 523310 638296 523316 638308
rect 523271 638268 523316 638296
rect 523310 638256 523316 638268
rect 523368 638256 523374 638308
rect 148042 638188 148048 638240
rect 148100 638228 148106 638240
rect 565078 638228 565084 638240
rect 148100 638200 565084 638228
rect 148100 638188 148106 638200
rect 565078 638188 565084 638200
rect 565136 638188 565142 638240
rect 126882 638120 126888 638172
rect 126940 638160 126946 638172
rect 544378 638160 544384 638172
rect 126940 638132 544384 638160
rect 126940 638120 126946 638132
rect 544378 638120 544384 638132
rect 544436 638120 544442 638172
rect 114462 638052 114468 638104
rect 114520 638092 114526 638104
rect 547138 638092 547144 638104
rect 114520 638064 547144 638092
rect 114520 638052 114526 638064
rect 547138 638052 547144 638064
rect 547196 638052 547202 638104
rect 102042 637984 102048 638036
rect 102100 638024 102106 638036
rect 548518 638024 548524 638036
rect 102100 637996 548524 638024
rect 102100 637984 102106 637996
rect 548518 637984 548524 637996
rect 548576 637984 548582 638036
rect 97902 637956 97908 637968
rect 97863 637928 97908 637956
rect 97902 637916 97908 637928
rect 97960 637916 97966 637968
rect 110322 637916 110328 637968
rect 110380 637956 110386 637968
rect 117133 637959 117191 637965
rect 117133 637956 117145 637959
rect 110380 637928 117145 637956
rect 110380 637916 110386 637928
rect 117133 637925 117145 637928
rect 117179 637925 117191 637959
rect 117133 637919 117191 637925
rect 122742 637916 122748 637968
rect 122800 637956 122806 637968
rect 576118 637956 576124 637968
rect 122800 637928 576124 637956
rect 122800 637916 122806 637928
rect 576118 637916 576124 637928
rect 576176 637916 576182 637968
rect 89530 637848 89536 637900
rect 89588 637888 89594 637900
rect 551278 637888 551284 637900
rect 89588 637860 551284 637888
rect 89588 637848 89594 637860
rect 551278 637848 551284 637860
rect 551336 637848 551342 637900
rect 117133 637823 117191 637829
rect 117133 637789 117145 637823
rect 117179 637820 117191 637823
rect 574738 637820 574744 637832
rect 117179 637792 574744 637820
rect 117179 637789 117191 637792
rect 117133 637783 117191 637789
rect 574738 637780 574744 637792
rect 574796 637780 574802 637832
rect 7558 637712 7564 637764
rect 7616 637752 7622 637764
rect 473357 637755 473415 637761
rect 473357 637752 473369 637755
rect 7616 637724 473369 637752
rect 7616 637712 7622 637724
rect 473357 637721 473369 637724
rect 473403 637721 473415 637755
rect 473357 637715 473415 637721
rect 97905 637687 97963 637693
rect 97905 637653 97917 637687
rect 97951 637684 97963 637687
rect 573358 637684 573364 637696
rect 97951 637656 573364 637684
rect 97951 637653 97963 637656
rect 97905 637647 97963 637653
rect 573358 637644 573364 637656
rect 573416 637644 573422 637696
rect 21358 637576 21364 637628
rect 21416 637616 21422 637628
rect 502521 637619 502579 637625
rect 502521 637616 502533 637619
rect 21416 637588 502533 637616
rect 21416 637576 21422 637588
rect 502521 637585 502533 637588
rect 502567 637585 502579 637619
rect 502521 637579 502579 637585
rect 35158 636828 35164 636880
rect 35216 636868 35222 636880
rect 523313 636871 523371 636877
rect 523313 636868 523325 636871
rect 35216 636840 523325 636868
rect 35216 636828 35222 636840
rect 523313 636837 523325 636840
rect 523359 636837 523371 636871
rect 523313 636831 523371 636837
rect 3326 632272 3332 632324
rect 3384 632312 3390 632324
rect 7650 632312 7656 632324
rect 3384 632284 7656 632312
rect 3384 632272 3390 632284
rect 7650 632272 7656 632284
rect 7708 632272 7714 632324
rect 530670 632000 530676 632052
rect 530728 632040 530734 632052
rect 579706 632040 579712 632052
rect 530728 632012 579712 632040
rect 530728 632000 530734 632012
rect 579706 632000 579712 632012
rect 579764 632000 579770 632052
rect 3602 619556 3608 619608
rect 3660 619596 3666 619608
rect 40862 619596 40868 619608
rect 3660 619568 40868 619596
rect 3660 619556 3666 619568
rect 40862 619556 40868 619568
rect 40920 619556 40926 619608
rect 538950 618196 538956 618248
rect 539008 618236 539014 618248
rect 579798 618236 579804 618248
rect 539008 618208 579804 618236
rect 539008 618196 539014 618208
rect 579798 618196 579804 618208
rect 579856 618196 579862 618248
rect 3050 607112 3056 607164
rect 3108 607152 3114 607164
rect 32490 607152 32496 607164
rect 3108 607124 32496 607152
rect 3108 607112 3114 607124
rect 32490 607112 32496 607124
rect 32548 607112 32554 607164
rect 565170 591948 565176 592000
rect 565228 591988 565234 592000
rect 580166 591988 580172 592000
rect 565228 591960 580172 591988
rect 565228 591948 565234 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 3326 580932 3332 580984
rect 3384 580972 3390 580984
rect 11790 580972 11796 580984
rect 3384 580944 11796 580972
rect 3384 580932 3390 580944
rect 11790 580932 11796 580944
rect 11848 580932 11854 580984
rect 569310 578144 569316 578196
rect 569368 578184 569374 578196
rect 580166 578184 580172 578196
rect 569368 578156 580172 578184
rect 569368 578144 569374 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 3326 567128 3332 567180
rect 3384 567168 3390 567180
rect 43530 567168 43536 567180
rect 3384 567140 43536 567168
rect 3384 567128 3390 567140
rect 43530 567128 43536 567140
rect 43588 567128 43594 567180
rect 537570 564340 537576 564392
rect 537628 564380 537634 564392
rect 580166 564380 580172 564392
rect 537628 564352 580172 564380
rect 537628 564340 537634 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3326 554684 3332 554736
rect 3384 554724 3390 554736
rect 33870 554724 33876 554736
rect 3384 554696 33876 554724
rect 3384 554684 3390 554696
rect 33870 554684 33876 554696
rect 33928 554684 33934 554736
rect 562410 538160 562416 538212
rect 562468 538200 562474 538212
rect 580166 538200 580172 538212
rect 562468 538172 580172 538200
rect 562468 538160 562474 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3326 528504 3332 528556
rect 3384 528544 3390 528556
rect 14550 528544 14556 528556
rect 3384 528516 14556 528544
rect 3384 528504 3390 528516
rect 14550 528504 14556 528516
rect 14608 528504 14614 528556
rect 558270 525716 558276 525768
rect 558328 525756 558334 525768
rect 580166 525756 580172 525768
rect 558328 525728 580172 525756
rect 558328 525716 558334 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 3142 516060 3148 516112
rect 3200 516100 3206 516112
rect 14458 516100 14464 516112
rect 3200 516072 14464 516100
rect 3200 516060 3206 516072
rect 14458 516060 14464 516072
rect 14516 516060 14522 516112
rect 536190 511912 536196 511964
rect 536248 511952 536254 511964
rect 580166 511952 580172 511964
rect 536248 511924 580172 511952
rect 536248 511912 536254 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 2958 502256 2964 502308
rect 3016 502296 3022 502308
rect 35250 502296 35256 502308
rect 3016 502268 35256 502296
rect 3016 502256 3022 502268
rect 35250 502256 35256 502268
rect 35308 502256 35314 502308
rect 561122 485732 561128 485784
rect 561180 485772 561186 485784
rect 580166 485772 580172 485784
rect 561180 485744 580172 485772
rect 561180 485732 561186 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3234 476008 3240 476060
rect 3292 476048 3298 476060
rect 15930 476048 15936 476060
rect 3292 476020 15936 476048
rect 3292 476008 3298 476020
rect 15930 476008 15936 476020
rect 15988 476008 15994 476060
rect 536098 471928 536104 471980
rect 536156 471968 536162 471980
rect 580166 471968 580172 471980
rect 536156 471940 580172 471968
rect 536156 471928 536162 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 3050 463632 3056 463684
rect 3108 463672 3114 463684
rect 15838 463672 15844 463684
rect 3108 463644 15844 463672
rect 3108 463632 3114 463644
rect 15838 463632 15844 463644
rect 15896 463632 15902 463684
rect 533430 458124 533436 458176
rect 533488 458164 533494 458176
rect 580166 458164 580172 458176
rect 533488 458136 580172 458164
rect 533488 458124 533494 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 40770 449868 40776 449880
rect 3384 449840 40776 449868
rect 3384 449828 3390 449840
rect 40770 449828 40776 449840
rect 40828 449828 40834 449880
rect 562318 431876 562324 431928
rect 562376 431916 562382 431928
rect 580166 431916 580172 431928
rect 562376 431888 580172 431916
rect 562376 431876 562382 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 17310 423620 17316 423632
rect 3384 423592 17316 423620
rect 3384 423580 3390 423592
rect 17310 423580 17316 423592
rect 17368 423580 17374 423632
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 17218 411244 17224 411256
rect 3016 411216 17224 411244
rect 3016 411204 3022 411216
rect 17218 411204 17224 411216
rect 17276 411204 17282 411256
rect 551370 405628 551376 405680
rect 551428 405668 551434 405680
rect 580166 405668 580172 405680
rect 551428 405640 580172 405668
rect 551428 405628 551434 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 50430 398800 50436 398812
rect 3384 398772 50436 398800
rect 3384 398760 3390 398772
rect 50430 398760 50436 398772
rect 50488 398760 50494 398812
rect 537478 379448 537484 379500
rect 537536 379488 537542 379500
rect 580166 379488 580172 379500
rect 537536 379460 580172 379488
rect 537536 379448 537542 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 372512 3332 372564
rect 3384 372552 3390 372564
rect 18690 372552 18696 372564
rect 3384 372524 18696 372552
rect 3384 372512 3390 372524
rect 18690 372512 18696 372524
rect 18748 372512 18754 372564
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 40678 358748 40684 358760
rect 3384 358720 40684 358748
rect 3384 358708 3390 358720
rect 40678 358708 40684 358720
rect 40736 358708 40742 358760
rect 548610 353200 548616 353252
rect 548668 353240 548674 353252
rect 580166 353240 580172 353252
rect 548668 353212 580172 353240
rect 548668 353200 548674 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 53190 346372 53196 346384
rect 3384 346344 53196 346372
rect 3384 346332 3390 346344
rect 53190 346332 53196 346344
rect 53248 346332 53254 346384
rect 565078 325592 565084 325644
rect 565136 325632 565142 325644
rect 579890 325632 579896 325644
rect 565136 325604 579896 325632
rect 565136 325592 565142 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 21450 320124 21456 320136
rect 3384 320096 21456 320124
rect 3384 320084 3390 320096
rect 21450 320084 21456 320096
rect 21508 320084 21514 320136
rect 532050 313216 532056 313268
rect 532108 313256 532114 313268
rect 580166 313256 580172 313268
rect 532108 313228 580172 313256
rect 532108 313216 532114 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 50338 306320 50344 306332
rect 3384 306292 50344 306320
rect 3384 306280 3390 306292
rect 50338 306280 50344 306292
rect 50396 306280 50402 306332
rect 547230 299412 547236 299464
rect 547288 299452 547294 299464
rect 579614 299452 579620 299464
rect 547288 299424 579620 299452
rect 547288 299412 547294 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 43438 293944 43444 293956
rect 3384 293916 43444 293944
rect 3384 293904 3390 293916
rect 43438 293904 43444 293916
rect 43496 293904 43502 293956
rect 538858 273164 538864 273216
rect 538916 273204 538922 273216
rect 579890 273204 579896 273216
rect 538916 273176 579896 273204
rect 538916 273164 538922 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 22738 267696 22744 267708
rect 3016 267668 22744 267696
rect 3016 267656 3022 267668
rect 22738 267656 22744 267668
rect 22796 267656 22802 267708
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 18598 255252 18604 255264
rect 3200 255224 18604 255252
rect 3200 255212 3206 255224
rect 18598 255212 18604 255224
rect 18656 255212 18662 255264
rect 544470 245556 544476 245608
rect 544528 245596 544534 245608
rect 580166 245596 580172 245608
rect 544528 245568 580172 245596
rect 544528 245556 544534 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 51718 241448 51724 241460
rect 3292 241420 51724 241448
rect 3292 241408 3298 241420
rect 51718 241408 51724 241420
rect 51776 241408 51782 241460
rect 576118 233180 576124 233232
rect 576176 233220 576182 233232
rect 579982 233220 579988 233232
rect 576176 233192 579988 233220
rect 576176 233180 576182 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 544378 219376 544384 219428
rect 544436 219416 544442 219428
rect 580166 219416 580172 219428
rect 544436 219388 580172 219416
rect 544436 219376 544442 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 25498 215268 25504 215280
rect 3384 215240 25504 215268
rect 3384 215228 3390 215240
rect 25498 215228 25504 215240
rect 25556 215228 25562 215280
rect 542998 206932 543004 206984
rect 543056 206972 543062 206984
rect 579798 206972 579804 206984
rect 543056 206944 579804 206972
rect 543056 206932 543062 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 574738 193128 574744 193180
rect 574796 193168 574802 193180
rect 580166 193168 580172 193180
rect 574796 193140 580172 193168
rect 574796 193128 574802 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3510 188844 3516 188896
rect 3568 188884 3574 188896
rect 7558 188884 7564 188896
rect 3568 188856 7564 188884
rect 3568 188844 3574 188856
rect 7558 188844 7564 188856
rect 7616 188844 7622 188896
rect 547138 179324 547144 179376
rect 547196 179364 547202 179376
rect 580166 179364 580172 179376
rect 547196 179336 580172 179364
rect 547196 179324 547202 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 531958 166948 531964 167000
rect 532016 166988 532022 167000
rect 580166 166988 580172 167000
rect 532016 166960 580172 166988
rect 532016 166948 532022 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 36538 164200 36544 164212
rect 3292 164172 36544 164200
rect 3292 164160 3298 164172
rect 36538 164160 36544 164172
rect 36596 164160 36602 164212
rect 573358 153144 573364 153196
rect 573416 153184 573422 153196
rect 580166 153184 580172 153196
rect 573416 153156 580172 153184
rect 573416 153144 573422 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 53098 150396 53104 150408
rect 3568 150368 53104 150396
rect 3568 150356 3574 150368
rect 53098 150356 53104 150368
rect 53156 150356 53162 150408
rect 548518 139340 548524 139392
rect 548576 139380 548582 139392
rect 580166 139380 580172 139392
rect 548576 139352 580172 139380
rect 548576 139340 548582 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 32398 137952 32404 137964
rect 3568 137924 32404 137952
rect 3568 137912 3574 137924
rect 32398 137912 32404 137924
rect 32456 137912 32462 137964
rect 530578 126896 530584 126948
rect 530636 126936 530642 126948
rect 580166 126936 580172 126948
rect 530636 126908 580172 126936
rect 530636 126896 530642 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 569218 113092 569224 113144
rect 569276 113132 569282 113144
rect 579798 113132 579804 113144
rect 569276 113104 579804 113132
rect 569276 113092 569282 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 39298 111772 39304 111784
rect 3200 111744 39304 111772
rect 3200 111732 3206 111744
rect 39298 111732 39304 111744
rect 39356 111732 39362 111784
rect 551278 100648 551284 100700
rect 551336 100688 551342 100700
rect 580166 100688 580172 100700
rect 551336 100660 580172 100688
rect 551336 100648 551342 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 21358 97968 21364 97980
rect 3568 97940 21364 97968
rect 3568 97928 3574 97940
rect 21358 97928 21364 97940
rect 21416 97928 21422 97980
rect 540238 86912 540244 86964
rect 540296 86952 540302 86964
rect 580166 86952 580172 86964
rect 540296 86924 580172 86952
rect 540296 86912 540302 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 11698 85524 11704 85536
rect 3568 85496 11704 85524
rect 3568 85484 3574 85496
rect 11698 85484 11704 85496
rect 11756 85484 11762 85536
rect 566458 73108 566464 73160
rect 566516 73148 566522 73160
rect 580166 73148 580172 73160
rect 566516 73120 580172 73148
rect 566516 73108 566522 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 47578 71720 47584 71732
rect 3568 71692 47584 71720
rect 3568 71680 3574 71692
rect 47578 71680 47584 71692
rect 47636 71680 47642 71732
rect 23382 63452 23388 63504
rect 23440 63492 23446 63504
rect 72602 63492 72608 63504
rect 23440 63464 72608 63492
rect 23440 63452 23446 63464
rect 72602 63452 72608 63464
rect 72660 63452 72666 63504
rect 84838 63452 84844 63504
rect 84896 63492 84902 63504
rect 102502 63492 102508 63504
rect 84896 63464 102508 63492
rect 84896 63452 84902 63464
rect 102502 63452 102508 63464
rect 102560 63452 102566 63504
rect 105538 63452 105544 63504
rect 105596 63492 105602 63504
rect 117038 63492 117044 63504
rect 105596 63464 117044 63492
rect 105596 63452 105602 63464
rect 117038 63452 117044 63464
rect 117096 63452 117102 63504
rect 119798 63452 119804 63504
rect 119856 63492 119862 63504
rect 150802 63492 150808 63504
rect 119856 63464 150808 63492
rect 119856 63452 119862 63464
rect 150802 63452 150808 63464
rect 150860 63452 150866 63504
rect 157242 63452 157248 63504
rect 157300 63492 157306 63504
rect 181714 63492 181720 63504
rect 157300 63464 181720 63492
rect 157300 63452 157306 63464
rect 181714 63452 181720 63464
rect 181772 63452 181778 63504
rect 183462 63452 183468 63504
rect 183520 63492 183526 63504
rect 202966 63492 202972 63504
rect 183520 63464 202972 63492
rect 183520 63452 183526 63464
rect 202966 63452 202972 63464
rect 203024 63452 203030 63504
rect 209682 63452 209688 63504
rect 209740 63492 209746 63504
rect 224218 63492 224224 63504
rect 209740 63464 224224 63492
rect 209740 63452 209746 63464
rect 224218 63452 224224 63464
rect 224276 63452 224282 63504
rect 229002 63452 229008 63504
rect 229060 63492 229066 63504
rect 240686 63492 240692 63504
rect 229060 63464 240692 63492
rect 229060 63452 229066 63464
rect 240686 63452 240692 63464
rect 240744 63452 240750 63504
rect 248322 63452 248328 63504
rect 248380 63492 248386 63504
rect 256142 63492 256148 63504
rect 248380 63464 256148 63492
rect 248380 63452 248386 63464
rect 256142 63452 256148 63464
rect 256200 63452 256206 63504
rect 499574 63452 499580 63504
rect 499632 63492 499638 63504
rect 538858 63492 538864 63504
rect 499632 63464 538864 63492
rect 499632 63452 499638 63464
rect 538858 63452 538864 63464
rect 538916 63452 538922 63504
rect 24762 63384 24768 63436
rect 24820 63424 24826 63436
rect 73522 63424 73528 63436
rect 24820 63396 73528 63424
rect 24820 63384 24826 63396
rect 73522 63384 73528 63396
rect 73580 63384 73586 63436
rect 87598 63384 87604 63436
rect 87656 63424 87662 63436
rect 105446 63424 105452 63436
rect 87656 63396 105452 63424
rect 87656 63384 87662 63396
rect 105446 63384 105452 63396
rect 105504 63384 105510 63436
rect 115842 63384 115848 63436
rect 115900 63424 115906 63436
rect 147950 63424 147956 63436
rect 115900 63396 147956 63424
rect 115900 63384 115906 63396
rect 147950 63384 147956 63396
rect 148008 63384 148014 63436
rect 153010 63384 153016 63436
rect 153068 63424 153074 63436
rect 177850 63424 177856 63436
rect 153068 63396 177856 63424
rect 153068 63384 153074 63396
rect 177850 63384 177856 63396
rect 177908 63384 177914 63436
rect 186222 63384 186228 63436
rect 186280 63424 186286 63436
rect 205910 63424 205916 63436
rect 186280 63396 205916 63424
rect 186280 63384 186286 63396
rect 205910 63384 205916 63396
rect 205968 63384 205974 63436
rect 211062 63384 211068 63436
rect 211120 63424 211126 63436
rect 225230 63424 225236 63436
rect 211120 63396 225236 63424
rect 211120 63384 211126 63396
rect 225230 63384 225236 63396
rect 225288 63384 225294 63436
rect 226242 63384 226248 63436
rect 226300 63424 226306 63436
rect 237742 63424 237748 63436
rect 226300 63396 237748 63424
rect 226300 63384 226306 63396
rect 237742 63384 237748 63396
rect 237800 63384 237806 63436
rect 240778 63384 240784 63436
rect 240836 63424 240842 63436
rect 249334 63424 249340 63436
rect 240836 63396 249340 63424
rect 240836 63384 240842 63396
rect 249334 63384 249340 63396
rect 249392 63384 249398 63436
rect 470594 63384 470600 63436
rect 470652 63424 470658 63436
rect 508498 63424 508504 63436
rect 470652 63396 508504 63424
rect 470652 63384 470658 63396
rect 508498 63384 508504 63396
rect 508556 63384 508562 63436
rect 509234 63384 509240 63436
rect 509292 63424 509298 63436
rect 548518 63424 548524 63436
rect 509292 63396 548524 63424
rect 509292 63384 509298 63396
rect 548518 63384 548524 63396
rect 548576 63384 548582 63436
rect 26142 63316 26148 63368
rect 26200 63356 26206 63368
rect 74534 63356 74540 63368
rect 26200 63328 74540 63356
rect 26200 63316 26206 63328
rect 74534 63316 74540 63328
rect 74592 63316 74598 63368
rect 75270 63316 75276 63368
rect 75328 63356 75334 63368
rect 99650 63356 99656 63368
rect 75328 63328 99656 63356
rect 75328 63316 75334 63328
rect 99650 63316 99656 63328
rect 99708 63316 99714 63368
rect 106182 63316 106188 63368
rect 106240 63356 106246 63368
rect 140222 63356 140228 63368
rect 106240 63328 140228 63356
rect 106240 63316 106246 63328
rect 140222 63316 140228 63328
rect 140280 63316 140286 63368
rect 148962 63316 148968 63368
rect 149020 63356 149026 63368
rect 174998 63356 175004 63368
rect 149020 63328 175004 63356
rect 149020 63316 149026 63328
rect 174998 63316 175004 63328
rect 175056 63316 175062 63368
rect 177942 63316 177948 63368
rect 178000 63356 178006 63368
rect 198182 63356 198188 63368
rect 178000 63328 198188 63356
rect 178000 63316 178006 63328
rect 198182 63316 198188 63328
rect 198240 63316 198246 63368
rect 198642 63316 198648 63368
rect 198700 63356 198706 63368
rect 215570 63356 215576 63368
rect 198700 63328 215576 63356
rect 198700 63316 198706 63328
rect 215570 63316 215576 63328
rect 215628 63316 215634 63368
rect 219250 63316 219256 63368
rect 219308 63356 219314 63368
rect 231946 63356 231952 63368
rect 219308 63328 231952 63356
rect 219308 63316 219314 63328
rect 231946 63316 231952 63328
rect 232004 63316 232010 63368
rect 233142 63316 233148 63368
rect 233200 63356 233206 63368
rect 243538 63356 243544 63368
rect 233200 63328 243544 63356
rect 233200 63316 233206 63328
rect 243538 63316 243544 63328
rect 243596 63316 243602 63368
rect 244182 63316 244188 63368
rect 244240 63356 244246 63368
rect 252278 63356 252284 63368
rect 244240 63328 252284 63356
rect 244240 63316 244246 63328
rect 252278 63316 252284 63328
rect 252336 63316 252342 63368
rect 334342 63316 334348 63368
rect 334400 63356 334406 63368
rect 335262 63356 335268 63368
rect 334400 63328 335268 63356
rect 334400 63316 334406 63328
rect 335262 63316 335268 63328
rect 335320 63316 335326 63368
rect 353662 63316 353668 63368
rect 353720 63356 353726 63368
rect 354582 63356 354588 63368
rect 353720 63328 354588 63356
rect 353720 63316 353726 63328
rect 354582 63316 354588 63328
rect 354640 63316 354646 63368
rect 372982 63316 372988 63368
rect 373040 63356 373046 63368
rect 373902 63356 373908 63368
rect 373040 63328 373908 63356
rect 373040 63316 373046 63328
rect 373902 63316 373908 63328
rect 373960 63316 373966 63368
rect 392302 63316 392308 63368
rect 392360 63356 392366 63368
rect 393222 63356 393228 63368
rect 392360 63328 393228 63356
rect 392360 63316 392366 63328
rect 393222 63316 393228 63328
rect 393280 63316 393286 63368
rect 411622 63316 411628 63368
rect 411680 63356 411686 63368
rect 412542 63356 412548 63368
rect 411680 63328 412548 63356
rect 411680 63316 411686 63328
rect 412542 63316 412548 63328
rect 412600 63316 412606 63368
rect 445478 63316 445484 63368
rect 445536 63356 445542 63368
rect 449158 63356 449164 63368
rect 445536 63328 449164 63356
rect 445536 63316 445542 63328
rect 449158 63316 449164 63328
rect 449216 63316 449222 63368
rect 457070 63316 457076 63368
rect 457128 63356 457134 63368
rect 471238 63356 471244 63368
rect 457128 63328 471244 63356
rect 457128 63316 457134 63328
rect 471238 63316 471244 63328
rect 471296 63316 471302 63368
rect 494698 63316 494704 63368
rect 494756 63356 494762 63368
rect 495342 63356 495348 63368
rect 494756 63328 495348 63356
rect 494756 63316 494762 63328
rect 495342 63316 495348 63328
rect 495400 63316 495406 63368
rect 533430 63356 533436 63368
rect 495452 63328 533436 63356
rect 20622 63248 20628 63300
rect 20680 63288 20686 63300
rect 69658 63288 69664 63300
rect 20680 63260 69664 63288
rect 20680 63248 20686 63260
rect 69658 63248 69664 63260
rect 69716 63248 69722 63300
rect 79410 63248 79416 63300
rect 79468 63288 79474 63300
rect 88058 63288 88064 63300
rect 79468 63260 88064 63288
rect 79468 63248 79474 63260
rect 88058 63248 88064 63260
rect 88116 63248 88122 63300
rect 90358 63248 90364 63300
rect 90416 63288 90422 63300
rect 97718 63288 97724 63300
rect 90416 63260 97724 63288
rect 90416 63248 90422 63260
rect 97718 63248 97724 63260
rect 97776 63248 97782 63300
rect 99282 63248 99288 63300
rect 99340 63288 99346 63300
rect 134426 63288 134432 63300
rect 99340 63260 134432 63288
rect 99340 63248 99346 63260
rect 134426 63248 134432 63260
rect 134484 63248 134490 63300
rect 138658 63248 138664 63300
rect 138716 63288 138722 63300
rect 152734 63288 152740 63300
rect 138716 63260 152740 63288
rect 138716 63248 138722 63260
rect 152734 63248 152740 63260
rect 152792 63248 152798 63300
rect 154482 63248 154488 63300
rect 154540 63288 154546 63300
rect 179782 63288 179788 63300
rect 154540 63260 179788 63288
rect 154540 63248 154546 63260
rect 179782 63248 179788 63260
rect 179840 63248 179846 63300
rect 180702 63248 180708 63300
rect 180760 63288 180766 63300
rect 201034 63288 201040 63300
rect 180760 63260 201040 63288
rect 180760 63248 180766 63260
rect 201034 63248 201040 63260
rect 201092 63248 201098 63300
rect 204162 63248 204168 63300
rect 204220 63288 204226 63300
rect 220354 63288 220360 63300
rect 204220 63260 220360 63288
rect 204220 63248 204226 63260
rect 220354 63248 220360 63260
rect 220412 63248 220418 63300
rect 223482 63248 223488 63300
rect 223540 63288 223546 63300
rect 235810 63288 235816 63300
rect 223540 63260 235816 63288
rect 223540 63248 223546 63260
rect 235810 63248 235816 63260
rect 235868 63248 235874 63300
rect 235902 63248 235908 63300
rect 235960 63288 235966 63300
rect 246482 63288 246488 63300
rect 235960 63260 246488 63288
rect 235960 63248 235966 63260
rect 246482 63248 246488 63260
rect 246540 63248 246546 63300
rect 454126 63248 454132 63300
rect 454184 63288 454190 63300
rect 468478 63288 468484 63300
rect 454184 63260 468484 63288
rect 454184 63248 454190 63260
rect 468478 63248 468484 63260
rect 468536 63248 468542 63300
rect 482186 63248 482192 63300
rect 482244 63288 482250 63300
rect 482922 63288 482928 63300
rect 482244 63260 482928 63288
rect 482244 63248 482250 63260
rect 482922 63248 482928 63260
rect 482980 63248 482986 63300
rect 493778 63248 493784 63300
rect 493836 63288 493842 63300
rect 495452 63288 495480 63328
rect 533430 63316 533436 63328
rect 533488 63316 533494 63368
rect 493836 63260 495480 63288
rect 493836 63248 493842 63260
rect 496630 63248 496636 63300
rect 496688 63288 496694 63300
rect 537478 63288 537484 63300
rect 496688 63260 537484 63288
rect 496688 63248 496694 63260
rect 537478 63248 537484 63260
rect 537536 63248 537542 63300
rect 10962 63180 10968 63232
rect 11020 63220 11026 63232
rect 61930 63220 61936 63232
rect 11020 63192 61936 63220
rect 11020 63180 11026 63192
rect 61930 63180 61936 63192
rect 61988 63180 61994 63232
rect 75089 63223 75147 63229
rect 75089 63189 75101 63223
rect 75135 63220 75147 63223
rect 77386 63220 77392 63232
rect 75135 63192 77392 63220
rect 75135 63189 75147 63192
rect 75089 63183 75147 63189
rect 77386 63180 77392 63192
rect 77444 63180 77450 63232
rect 77938 63180 77944 63232
rect 77996 63220 78002 63232
rect 88978 63220 88984 63232
rect 77996 63192 88984 63220
rect 77996 63180 78002 63192
rect 88978 63180 88984 63192
rect 89036 63180 89042 63232
rect 93762 63180 93768 63232
rect 93820 63220 93826 63232
rect 129550 63220 129556 63232
rect 93820 63192 129556 63220
rect 93820 63180 93826 63192
rect 129550 63180 129556 63192
rect 129608 63180 129614 63232
rect 134518 63180 134524 63232
rect 134576 63220 134582 63232
rect 144086 63220 144092 63232
rect 134576 63192 144092 63220
rect 134576 63180 134582 63192
rect 144086 63180 144092 63192
rect 144144 63180 144150 63232
rect 144822 63180 144828 63232
rect 144880 63220 144886 63232
rect 172054 63220 172060 63232
rect 144880 63192 172060 63220
rect 144880 63180 144886 63192
rect 172054 63180 172060 63192
rect 172112 63180 172118 63232
rect 175182 63180 175188 63232
rect 175240 63220 175246 63232
rect 196250 63220 196256 63232
rect 175240 63192 196256 63220
rect 175240 63180 175246 63192
rect 196250 63180 196256 63192
rect 196308 63180 196314 63232
rect 197262 63180 197268 63232
rect 197320 63220 197326 63232
rect 214558 63220 214564 63232
rect 197320 63192 214564 63220
rect 197320 63180 197326 63192
rect 214558 63180 214564 63192
rect 214616 63180 214622 63232
rect 215202 63180 215208 63232
rect 215260 63220 215266 63232
rect 229094 63220 229100 63232
rect 215260 63192 229100 63220
rect 215260 63180 215266 63192
rect 229094 63180 229100 63192
rect 229152 63180 229158 63232
rect 231762 63180 231768 63232
rect 231820 63220 231826 63232
rect 242618 63220 242624 63232
rect 231820 63192 242624 63220
rect 231820 63180 231826 63192
rect 242618 63180 242624 63192
rect 242676 63180 242682 63232
rect 246942 63180 246948 63232
rect 247000 63220 247006 63232
rect 255130 63220 255136 63232
rect 247000 63192 255136 63220
rect 247000 63180 247006 63192
rect 255130 63180 255136 63192
rect 255188 63180 255194 63232
rect 439682 63180 439688 63232
rect 439740 63220 439746 63232
rect 440142 63220 440148 63232
rect 439740 63192 440148 63220
rect 439740 63180 439746 63192
rect 440142 63180 440148 63192
rect 440200 63180 440206 63232
rect 462866 63180 462872 63232
rect 462924 63220 462930 63232
rect 482278 63220 482284 63232
rect 462924 63192 482284 63220
rect 462924 63180 462930 63192
rect 482278 63180 482284 63192
rect 482336 63180 482342 63232
rect 489914 63180 489920 63232
rect 489972 63220 489978 63232
rect 497553 63223 497611 63229
rect 497553 63220 497565 63223
rect 489972 63192 497565 63220
rect 489972 63180 489978 63192
rect 497553 63189 497565 63192
rect 497599 63189 497611 63223
rect 497553 63183 497611 63189
rect 506290 63180 506296 63232
rect 506348 63220 506354 63232
rect 547138 63220 547144 63232
rect 506348 63192 547144 63220
rect 506348 63180 506354 63192
rect 547138 63180 547144 63192
rect 547196 63180 547202 63232
rect 12342 63112 12348 63164
rect 12400 63152 12406 63164
rect 62942 63152 62948 63164
rect 12400 63124 62948 63152
rect 12400 63112 12406 63124
rect 62942 63112 62948 63124
rect 63000 63112 63006 63164
rect 64138 63112 64144 63164
rect 64196 63152 64202 63164
rect 83182 63152 83188 63164
rect 64196 63124 83188 63152
rect 64196 63112 64202 63124
rect 83182 63112 83188 63124
rect 83240 63112 83246 63164
rect 86862 63112 86868 63164
rect 86920 63152 86926 63164
rect 123754 63152 123760 63164
rect 86920 63124 123760 63152
rect 86920 63112 86926 63124
rect 123754 63112 123760 63124
rect 123812 63112 123818 63164
rect 124122 63112 124128 63164
rect 124180 63152 124186 63164
rect 154666 63152 154672 63164
rect 124180 63124 154672 63152
rect 124180 63112 124186 63124
rect 154666 63112 154672 63124
rect 154724 63112 154730 63164
rect 155862 63112 155868 63164
rect 155920 63152 155926 63164
rect 180794 63152 180800 63164
rect 155920 63124 180800 63152
rect 155920 63112 155926 63124
rect 180794 63112 180800 63124
rect 180852 63112 180858 63164
rect 182082 63112 182088 63164
rect 182140 63152 182146 63164
rect 202046 63152 202052 63164
rect 182140 63124 202052 63152
rect 182140 63112 182146 63124
rect 202046 63112 202052 63124
rect 202104 63112 202110 63164
rect 205542 63112 205548 63164
rect 205600 63152 205606 63164
rect 221366 63152 221372 63164
rect 205600 63124 221372 63152
rect 205600 63112 205606 63124
rect 221366 63112 221372 63124
rect 221424 63112 221430 63164
rect 222102 63112 222108 63164
rect 222160 63152 222166 63164
rect 234890 63152 234896 63164
rect 222160 63124 234896 63152
rect 222160 63112 222166 63124
rect 234890 63112 234896 63124
rect 234948 63112 234954 63164
rect 237282 63112 237288 63164
rect 237340 63152 237346 63164
rect 247402 63152 247408 63164
rect 237340 63124 247408 63152
rect 237340 63112 237346 63124
rect 247402 63112 247408 63124
rect 247460 63112 247466 63164
rect 255958 63112 255964 63164
rect 256016 63152 256022 63164
rect 261938 63152 261944 63164
rect 256016 63124 261944 63152
rect 256016 63112 256022 63124
rect 261938 63112 261944 63124
rect 261996 63112 262002 63164
rect 328546 63112 328552 63164
rect 328604 63152 328610 63164
rect 329650 63152 329656 63164
rect 328604 63124 329656 63152
rect 328604 63112 328610 63124
rect 329650 63112 329656 63124
rect 329708 63112 329714 63164
rect 367186 63112 367192 63164
rect 367244 63152 367250 63164
rect 368290 63152 368296 63164
rect 367244 63124 368296 63152
rect 367244 63112 367250 63124
rect 368290 63112 368296 63124
rect 368348 63112 368354 63164
rect 386506 63112 386512 63164
rect 386564 63152 386570 63164
rect 387610 63152 387616 63164
rect 386564 63124 387616 63152
rect 386564 63112 386570 63124
rect 387610 63112 387616 63124
rect 387668 63112 387674 63164
rect 405826 63112 405832 63164
rect 405884 63152 405890 63164
rect 406930 63152 406936 63164
rect 405884 63124 406936 63152
rect 405884 63112 405890 63124
rect 406930 63112 406936 63124
rect 406988 63112 406994 63164
rect 440602 63112 440608 63164
rect 440660 63152 440666 63164
rect 441522 63152 441528 63164
rect 440660 63124 441528 63152
rect 440660 63112 440666 63124
rect 441522 63112 441528 63124
rect 441580 63112 441586 63164
rect 451274 63112 451280 63164
rect 451332 63152 451338 63164
rect 467098 63152 467104 63164
rect 451332 63124 467104 63152
rect 451332 63112 451338 63124
rect 467098 63112 467104 63124
rect 467156 63112 467162 63164
rect 467650 63112 467656 63164
rect 467708 63152 467714 63164
rect 502978 63152 502984 63164
rect 467708 63124 502984 63152
rect 467708 63112 467714 63124
rect 502978 63112 502984 63124
rect 503036 63112 503042 63164
rect 503438 63112 503444 63164
rect 503496 63152 503502 63164
rect 544378 63152 544384 63164
rect 503496 63124 544384 63152
rect 503496 63112 503502 63124
rect 544378 63112 544384 63124
rect 544436 63112 544442 63164
rect 65518 63044 65524 63096
rect 65576 63084 65582 63096
rect 89990 63084 89996 63096
rect 65576 63056 89996 63084
rect 65576 63044 65582 63056
rect 89990 63044 89996 63056
rect 90048 63044 90054 63096
rect 95142 63044 95148 63096
rect 95200 63084 95206 63096
rect 131482 63084 131488 63096
rect 95200 63056 131488 63084
rect 95200 63044 95206 63056
rect 131482 63044 131488 63056
rect 131540 63044 131546 63096
rect 142062 63044 142068 63096
rect 142120 63084 142126 63096
rect 169202 63084 169208 63096
rect 142120 63056 169208 63084
rect 142120 63044 142126 63056
rect 169202 63044 169208 63056
rect 169260 63044 169266 63096
rect 169662 63044 169668 63096
rect 169720 63084 169726 63096
rect 192386 63084 192392 63096
rect 169720 63056 192392 63084
rect 169720 63044 169726 63056
rect 192386 63044 192392 63056
rect 192444 63044 192450 63096
rect 194410 63044 194416 63096
rect 194468 63084 194474 63096
rect 211706 63084 211712 63096
rect 194468 63056 211712 63084
rect 194468 63044 194474 63056
rect 211706 63044 211712 63056
rect 211764 63044 211770 63096
rect 212442 63044 212448 63096
rect 212500 63084 212506 63096
rect 227162 63084 227168 63096
rect 212500 63056 227168 63084
rect 212500 63044 212506 63056
rect 227162 63044 227168 63056
rect 227220 63044 227226 63096
rect 227622 63044 227628 63096
rect 227680 63084 227686 63096
rect 239674 63084 239680 63096
rect 227680 63056 239680 63084
rect 227680 63044 227686 63056
rect 239674 63044 239680 63056
rect 239732 63044 239738 63096
rect 241422 63044 241428 63096
rect 241480 63084 241486 63096
rect 250346 63084 250352 63096
rect 241480 63056 250352 63084
rect 241480 63044 241486 63056
rect 250346 63044 250352 63056
rect 250404 63044 250410 63096
rect 251082 63044 251088 63096
rect 251140 63084 251146 63096
rect 258074 63084 258080 63096
rect 251140 63056 258080 63084
rect 251140 63044 251146 63056
rect 258074 63044 258080 63056
rect 258132 63044 258138 63096
rect 267642 63044 267648 63096
rect 267700 63084 267706 63096
rect 271598 63084 271604 63096
rect 267700 63056 271604 63084
rect 267700 63044 267706 63056
rect 271598 63044 271604 63056
rect 271656 63044 271662 63096
rect 422294 63044 422300 63096
rect 422352 63084 422358 63096
rect 436646 63084 436652 63096
rect 422352 63056 436652 63084
rect 422352 63044 422358 63056
rect 436646 63044 436652 63056
rect 436704 63044 436710 63096
rect 444466 63044 444472 63096
rect 444524 63084 444530 63096
rect 464338 63084 464344 63096
rect 444524 63056 464344 63084
rect 444524 63044 444530 63056
rect 464338 63044 464344 63056
rect 464396 63044 464402 63096
rect 474458 63044 474464 63096
rect 474516 63084 474522 63096
rect 490558 63084 490564 63096
rect 474516 63056 490564 63084
rect 474516 63044 474522 63056
rect 490558 63044 490564 63056
rect 490616 63044 490622 63096
rect 490834 63044 490840 63096
rect 490892 63084 490898 63096
rect 532050 63084 532056 63096
rect 490892 63056 532056 63084
rect 490892 63044 490898 63056
rect 532050 63044 532056 63056
rect 532108 63044 532114 63096
rect 16482 62976 16488 63028
rect 16540 63016 16546 63028
rect 66806 63016 66812 63028
rect 16540 62988 66812 63016
rect 16540 62976 16546 62988
rect 66806 62976 66812 62988
rect 66864 62976 66870 63028
rect 72418 62976 72424 63028
rect 72476 63016 72482 63028
rect 78398 63016 78404 63028
rect 72476 62988 78404 63016
rect 72476 62976 72482 62988
rect 78398 62976 78404 62988
rect 78456 62976 78462 63028
rect 78493 63019 78551 63025
rect 78493 62985 78505 63019
rect 78539 63016 78551 63019
rect 78539 62988 79456 63016
rect 78539 62985 78551 62988
rect 78493 62979 78551 62985
rect 13722 62908 13728 62960
rect 13780 62948 13786 62960
rect 64874 62948 64880 62960
rect 13780 62920 64880 62948
rect 13780 62908 13786 62920
rect 64874 62908 64880 62920
rect 64932 62908 64938 62960
rect 71682 62908 71688 62960
rect 71740 62948 71746 62960
rect 79428 62948 79456 62988
rect 81342 62976 81348 63028
rect 81400 63016 81406 63028
rect 119890 63016 119896 63028
rect 81400 62988 119896 63016
rect 81400 62976 81406 62988
rect 119890 62976 119896 62988
rect 119948 62976 119954 63028
rect 119982 62976 119988 63028
rect 120040 63016 120046 63028
rect 151814 63016 151820 63028
rect 120040 62988 151820 63016
rect 120040 62976 120046 62988
rect 151814 62976 151820 62988
rect 151872 62976 151878 63028
rect 153102 62976 153108 63028
rect 153160 63016 153166 63028
rect 178862 63016 178868 63028
rect 153160 62988 178868 63016
rect 153160 62976 153166 62988
rect 178862 62976 178868 62988
rect 178920 62976 178926 63028
rect 179322 62976 179328 63028
rect 179380 63016 179386 63028
rect 200114 63016 200120 63028
rect 179380 62988 200120 63016
rect 179380 62976 179386 62988
rect 200114 62976 200120 62988
rect 200172 62976 200178 63028
rect 206922 62976 206928 63028
rect 206980 63016 206986 63028
rect 222286 63016 222292 63028
rect 206980 62988 222292 63016
rect 206980 62976 206986 62988
rect 222286 62976 222292 62988
rect 222344 62976 222350 63028
rect 224862 62976 224868 63028
rect 224920 63016 224926 63028
rect 236822 63016 236828 63028
rect 224920 62988 236828 63016
rect 224920 62976 224926 62988
rect 236822 62976 236828 62988
rect 236880 62976 236886 63028
rect 238662 62976 238668 63028
rect 238720 63016 238726 63028
rect 248414 63016 248420 63028
rect 238720 62988 248420 63016
rect 238720 62976 238726 62988
rect 248414 62976 248420 62988
rect 248472 62976 248478 63028
rect 257982 62976 257988 63028
rect 258040 63016 258046 63028
rect 263870 63016 263876 63028
rect 258040 62988 263876 63016
rect 258040 62976 258046 62988
rect 263870 62976 263876 62988
rect 263928 62976 263934 63028
rect 311158 62976 311164 63028
rect 311216 63016 311222 63028
rect 311802 63016 311808 63028
rect 311216 62988 311808 63016
rect 311216 62976 311222 62988
rect 311802 62976 311808 62988
rect 311860 62976 311866 63028
rect 318886 62976 318892 63028
rect 318944 63016 318950 63028
rect 321002 63016 321008 63028
rect 318944 62988 321008 63016
rect 318944 62976 318950 62988
rect 321002 62976 321008 62988
rect 321060 62976 321066 63028
rect 330478 62976 330484 63028
rect 330536 63016 330542 63028
rect 331122 63016 331128 63028
rect 330536 62988 331128 63016
rect 330536 62976 330542 62988
rect 331122 62976 331128 62988
rect 331180 62976 331186 63028
rect 349798 62976 349804 63028
rect 349856 63016 349862 63028
rect 350442 63016 350448 63028
rect 349856 62988 350448 63016
rect 349856 62976 349862 62988
rect 350442 62976 350448 62988
rect 350500 62976 350506 63028
rect 369118 62976 369124 63028
rect 369176 63016 369182 63028
rect 369762 63016 369768 63028
rect 369176 62988 369768 63016
rect 369176 62976 369182 62988
rect 369762 62976 369768 62988
rect 369820 62976 369826 63028
rect 388438 62976 388444 63028
rect 388496 63016 388502 63028
rect 389082 63016 389088 63028
rect 388496 62988 389088 63016
rect 388496 62976 388502 62988
rect 389082 62976 389088 62988
rect 389140 62976 389146 63028
rect 407758 62976 407764 63028
rect 407816 63016 407822 63028
rect 408402 63016 408408 63028
rect 407816 62988 408408 63016
rect 407816 62976 407822 62988
rect 408402 62976 408408 62988
rect 408460 62976 408466 63028
rect 421282 62976 421288 63028
rect 421340 63016 421346 63028
rect 422202 63016 422208 63028
rect 421340 62988 422208 63016
rect 421340 62976 421346 62988
rect 422202 62976 422208 62988
rect 422260 62976 422266 63028
rect 427078 62976 427084 63028
rect 427136 63016 427142 63028
rect 427722 63016 427728 63028
rect 427136 62988 427728 63016
rect 427136 62976 427142 62988
rect 427722 62976 427728 62988
rect 427780 62976 427786 63028
rect 437750 62976 437756 63028
rect 437808 63016 437814 63028
rect 454678 63016 454684 63028
rect 437808 62988 454684 63016
rect 437808 62976 437814 62988
rect 454678 62976 454684 62988
rect 454736 62976 454742 63028
rect 463786 62976 463792 63028
rect 463844 63016 463850 63028
rect 500310 63016 500316 63028
rect 463844 62988 500316 63016
rect 463844 62976 463850 62988
rect 500310 62976 500316 62988
rect 500368 62976 500374 63028
rect 500494 62976 500500 63028
rect 500552 63016 500558 63028
rect 542998 63016 543004 63028
rect 500552 62988 543004 63016
rect 500552 62976 500558 62988
rect 542998 62976 543004 62988
rect 543056 62976 543062 63028
rect 85114 62948 85120 62960
rect 71740 62920 79364 62948
rect 79428 62920 85120 62948
rect 71740 62908 71746 62920
rect 6822 62840 6828 62892
rect 6880 62880 6886 62892
rect 59078 62880 59084 62892
rect 6880 62852 59084 62880
rect 6880 62840 6886 62852
rect 59078 62840 59084 62852
rect 59136 62840 59142 62892
rect 62758 62840 62764 62892
rect 62816 62880 62822 62892
rect 70670 62880 70676 62892
rect 62816 62852 70676 62880
rect 62816 62840 62822 62852
rect 70670 62840 70676 62852
rect 70728 62840 70734 62892
rect 73798 62840 73804 62892
rect 73856 62880 73862 62892
rect 76466 62880 76472 62892
rect 73856 62852 76472 62880
rect 73856 62840 73862 62852
rect 76466 62840 76472 62852
rect 76524 62840 76530 62892
rect 76558 62840 76564 62892
rect 76616 62880 76622 62892
rect 78493 62883 78551 62889
rect 78493 62880 78505 62883
rect 76616 62852 78505 62880
rect 76616 62840 76622 62852
rect 78493 62849 78505 62852
rect 78539 62849 78551 62883
rect 79336 62880 79364 62920
rect 85114 62908 85120 62920
rect 85172 62908 85178 62960
rect 88242 62908 88248 62960
rect 88300 62948 88306 62960
rect 125686 62948 125692 62960
rect 88300 62920 125692 62948
rect 88300 62908 88306 62920
rect 125686 62908 125692 62920
rect 125744 62908 125750 62960
rect 128998 62908 129004 62960
rect 129056 62948 129062 62960
rect 138290 62948 138296 62960
rect 129056 62920 138296 62948
rect 129056 62908 129062 62920
rect 138290 62908 138296 62920
rect 138348 62908 138354 62960
rect 143442 62908 143448 62960
rect 143500 62948 143506 62960
rect 170122 62948 170128 62960
rect 143500 62920 170128 62948
rect 143500 62908 143506 62920
rect 170122 62908 170128 62920
rect 170180 62908 170186 62960
rect 171042 62908 171048 62960
rect 171100 62948 171106 62960
rect 193306 62948 193312 62960
rect 171100 62920 193312 62948
rect 171100 62908 171106 62920
rect 193306 62908 193312 62920
rect 193364 62908 193370 62960
rect 194502 62908 194508 62960
rect 194560 62948 194566 62960
rect 212626 62948 212632 62960
rect 194560 62920 212632 62948
rect 194560 62908 194566 62920
rect 212626 62908 212632 62920
rect 212684 62908 212690 62960
rect 213822 62908 213828 62960
rect 213880 62948 213886 62960
rect 228082 62948 228088 62960
rect 213880 62920 228088 62948
rect 213880 62908 213886 62920
rect 228082 62908 228088 62920
rect 228140 62908 228146 62960
rect 230382 62908 230388 62960
rect 230440 62948 230446 62960
rect 241606 62948 241612 62960
rect 230440 62920 241612 62948
rect 230440 62908 230446 62920
rect 241606 62908 241612 62920
rect 241664 62908 241670 62960
rect 242802 62908 242808 62960
rect 242860 62948 242866 62960
rect 251266 62948 251272 62960
rect 242860 62920 251272 62948
rect 242860 62908 242866 62920
rect 251266 62908 251272 62920
rect 251324 62908 251330 62960
rect 266998 62908 267004 62960
rect 267056 62948 267062 62960
rect 270586 62948 270592 62960
rect 267056 62920 270592 62948
rect 267056 62908 267062 62920
rect 270586 62908 270592 62920
rect 270644 62908 270650 62960
rect 423214 62908 423220 62960
rect 423272 62948 423278 62960
rect 423272 62920 431954 62948
rect 423272 62908 423278 62920
rect 112162 62880 112168 62892
rect 79336 62852 112168 62880
rect 78493 62843 78551 62849
rect 112162 62840 112168 62852
rect 112220 62840 112226 62892
rect 113082 62840 113088 62892
rect 113140 62880 113146 62892
rect 146018 62880 146024 62892
rect 113140 62852 146024 62880
rect 113140 62840 113146 62852
rect 146018 62840 146024 62852
rect 146076 62840 146082 62892
rect 150342 62840 150348 62892
rect 150400 62880 150406 62892
rect 175918 62880 175924 62892
rect 150400 62852 175924 62880
rect 150400 62840 150406 62852
rect 175918 62840 175924 62852
rect 175976 62840 175982 62892
rect 177850 62840 177856 62892
rect 177908 62880 177914 62892
rect 199102 62880 199108 62892
rect 177908 62852 199108 62880
rect 177908 62840 177914 62852
rect 199102 62840 199108 62852
rect 199160 62840 199166 62892
rect 202690 62840 202696 62892
rect 202748 62880 202754 62892
rect 219434 62880 219440 62892
rect 202748 62852 219440 62880
rect 202748 62840 202754 62852
rect 219434 62840 219440 62852
rect 219492 62840 219498 62892
rect 220722 62840 220728 62892
rect 220780 62880 220786 62892
rect 233878 62880 233884 62892
rect 220780 62852 233884 62880
rect 220780 62840 220786 62852
rect 233878 62840 233884 62852
rect 233936 62840 233942 62892
rect 234522 62840 234528 62892
rect 234580 62880 234586 62892
rect 244550 62880 244556 62892
rect 234580 62852 244556 62880
rect 234580 62840 234586 62852
rect 244550 62840 244556 62852
rect 244608 62840 244614 62892
rect 245562 62840 245568 62892
rect 245620 62880 245626 62892
rect 254210 62880 254216 62892
rect 245620 62852 254216 62880
rect 245620 62840 245626 62852
rect 254210 62840 254216 62852
rect 254268 62840 254274 62892
rect 256602 62840 256608 62892
rect 256660 62880 256666 62892
rect 262858 62880 262864 62892
rect 256660 62852 262864 62880
rect 256660 62840 256666 62852
rect 262858 62840 262864 62852
rect 262916 62840 262922 62892
rect 327626 62840 327632 62892
rect 327684 62880 327690 62892
rect 328362 62880 328368 62892
rect 327684 62852 328368 62880
rect 327684 62840 327690 62852
rect 328362 62840 328368 62852
rect 328420 62840 328426 62892
rect 346946 62840 346952 62892
rect 347004 62880 347010 62892
rect 347682 62880 347688 62892
rect 347004 62852 347688 62880
rect 347004 62840 347010 62852
rect 347682 62840 347688 62852
rect 347740 62840 347746 62892
rect 366266 62840 366272 62892
rect 366324 62880 366330 62892
rect 367002 62880 367008 62892
rect 366324 62852 367008 62880
rect 366324 62840 366330 62852
rect 367002 62840 367008 62852
rect 367060 62840 367066 62892
rect 385586 62840 385592 62892
rect 385644 62880 385650 62892
rect 386322 62880 386328 62892
rect 385644 62852 386328 62880
rect 385644 62840 385650 62852
rect 386322 62840 386328 62852
rect 386380 62840 386386 62892
rect 404906 62840 404912 62892
rect 404964 62880 404970 62892
rect 405642 62880 405648 62892
rect 404964 62852 405648 62880
rect 404964 62840 404970 62852
rect 405642 62840 405648 62852
rect 405700 62840 405706 62892
rect 416498 62840 416504 62892
rect 416556 62880 416562 62892
rect 416556 62852 422294 62880
rect 416556 62840 416562 62852
rect 4062 62772 4068 62824
rect 4120 62812 4126 62824
rect 57146 62812 57152 62824
rect 4120 62784 57152 62812
rect 4120 62772 4126 62784
rect 57146 62772 57152 62784
rect 57204 62772 57210 62824
rect 57882 62772 57888 62824
rect 57940 62812 57946 62824
rect 100570 62812 100576 62824
rect 57940 62784 100576 62812
rect 57940 62772 57946 62784
rect 100570 62772 100576 62784
rect 100628 62772 100634 62824
rect 103422 62772 103428 62824
rect 103480 62812 103486 62824
rect 137278 62812 137284 62824
rect 103480 62784 137284 62812
rect 103480 62772 103486 62784
rect 137278 62772 137284 62784
rect 137336 62772 137342 62824
rect 139302 62772 139308 62824
rect 139360 62812 139366 62824
rect 167270 62812 167276 62824
rect 139360 62784 167276 62812
rect 139360 62772 139366 62784
rect 167270 62772 167276 62784
rect 167328 62772 167334 62824
rect 168282 62772 168288 62824
rect 168340 62812 168346 62824
rect 190454 62812 190460 62824
rect 168340 62784 190460 62812
rect 168340 62772 168346 62784
rect 190454 62772 190460 62784
rect 190512 62772 190518 62824
rect 191742 62772 191748 62824
rect 191800 62812 191806 62824
rect 209774 62812 209780 62824
rect 191800 62784 209780 62812
rect 191800 62772 191806 62784
rect 209774 62772 209780 62784
rect 209832 62772 209838 62824
rect 210970 62772 210976 62824
rect 211028 62812 211034 62824
rect 226150 62812 226156 62824
rect 211028 62784 226156 62812
rect 211028 62772 211034 62784
rect 226150 62772 226156 62784
rect 226208 62772 226214 62824
rect 227530 62772 227536 62824
rect 227588 62812 227594 62824
rect 238754 62812 238760 62824
rect 227588 62784 238760 62812
rect 227588 62772 227594 62784
rect 238754 62772 238760 62784
rect 238812 62772 238818 62824
rect 244090 62772 244096 62824
rect 244148 62812 244154 62824
rect 253198 62812 253204 62824
rect 244148 62784 253204 62812
rect 244148 62772 244154 62784
rect 253198 62772 253204 62784
rect 253256 62772 253262 62824
rect 253842 62772 253848 62824
rect 253900 62812 253906 62824
rect 260926 62812 260932 62824
rect 253900 62784 260932 62812
rect 253900 62772 253906 62784
rect 260926 62772 260932 62784
rect 260984 62772 260990 62824
rect 277210 62772 277216 62824
rect 277268 62812 277274 62824
rect 280246 62812 280252 62824
rect 277268 62784 280252 62812
rect 277268 62772 277274 62784
rect 280246 62772 280252 62784
rect 280304 62772 280310 62824
rect 340138 62772 340144 62824
rect 340196 62812 340202 62824
rect 340782 62812 340788 62824
rect 340196 62784 340788 62812
rect 340196 62772 340202 62784
rect 340782 62772 340788 62784
rect 340840 62772 340846 62824
rect 359458 62772 359464 62824
rect 359516 62812 359522 62824
rect 360102 62812 360108 62824
rect 359516 62784 360108 62812
rect 359516 62772 359522 62784
rect 360102 62772 360108 62784
rect 360160 62772 360166 62824
rect 378778 62772 378784 62824
rect 378836 62812 378842 62824
rect 379422 62812 379428 62824
rect 378836 62784 379428 62812
rect 378836 62772 378842 62784
rect 379422 62772 379428 62784
rect 379480 62772 379486 62824
rect 398098 62772 398104 62824
rect 398156 62812 398162 62824
rect 398742 62812 398748 62824
rect 398156 62784 398748 62812
rect 398156 62772 398162 62784
rect 398742 62772 398748 62784
rect 398800 62772 398806 62824
rect 417418 62772 417424 62824
rect 417476 62812 417482 62824
rect 418062 62812 418068 62824
rect 417476 62784 418068 62812
rect 417476 62772 417482 62784
rect 418062 62772 418068 62784
rect 418120 62772 418126 62824
rect 422266 62812 422294 62852
rect 424226 62840 424232 62892
rect 424284 62880 424290 62892
rect 424962 62880 424968 62892
rect 424284 62852 424968 62880
rect 424284 62840 424290 62852
rect 424962 62840 424968 62852
rect 425020 62840 425026 62892
rect 431926 62880 431954 62920
rect 434806 62908 434812 62960
rect 434864 62948 434870 62960
rect 465166 62948 465172 62960
rect 434864 62920 465172 62948
rect 434864 62908 434870 62920
rect 465166 62908 465172 62920
rect 465224 62908 465230 62960
rect 468662 62908 468668 62960
rect 468720 62948 468726 62960
rect 487798 62948 487804 62960
rect 468720 62920 487804 62948
rect 468720 62908 468726 62920
rect 487798 62908 487804 62920
rect 487856 62908 487862 62960
rect 491846 62908 491852 62960
rect 491904 62948 491910 62960
rect 535454 62948 535460 62960
rect 491904 62920 535460 62948
rect 491904 62908 491910 62920
rect 535454 62908 535460 62920
rect 535512 62908 535518 62960
rect 446306 62880 446312 62892
rect 431926 62852 446312 62880
rect 446306 62840 446312 62852
rect 446364 62840 446370 62892
rect 464798 62840 464804 62892
rect 464856 62880 464862 62892
rect 464856 62852 489914 62880
rect 464856 62840 464862 62852
rect 431218 62812 431224 62824
rect 422266 62784 431224 62812
rect 431218 62772 431224 62784
rect 431276 62772 431282 62824
rect 442534 62772 442540 62824
rect 442592 62812 442598 62824
rect 473998 62812 474004 62824
rect 442592 62784 474004 62812
rect 442592 62772 442598 62784
rect 473998 62772 474004 62784
rect 474056 62772 474062 62824
rect 489886 62812 489914 62852
rect 492766 62840 492772 62892
rect 492824 62880 492830 62892
rect 493962 62880 493968 62892
rect 492824 62852 493968 62880
rect 492824 62840 492830 62852
rect 493962 62840 493968 62852
rect 494020 62840 494026 62892
rect 497642 62840 497648 62892
rect 497700 62880 497706 62892
rect 541618 62880 541624 62892
rect 497700 62852 541624 62880
rect 497700 62840 497706 62852
rect 541618 62840 541624 62852
rect 541676 62840 541682 62892
rect 497458 62812 497464 62824
rect 489886 62784 497464 62812
rect 497458 62772 497464 62784
rect 497516 62772 497522 62824
rect 497553 62815 497611 62821
rect 497553 62781 497565 62815
rect 497599 62812 497611 62815
rect 529198 62812 529204 62824
rect 497599 62784 529204 62812
rect 497599 62781 497611 62784
rect 497553 62775 497611 62781
rect 529198 62772 529204 62784
rect 529256 62772 529262 62824
rect 529474 62772 529480 62824
rect 529532 62812 529538 62824
rect 582377 62815 582435 62821
rect 582377 62812 582389 62815
rect 529532 62784 582389 62812
rect 529532 62772 529538 62784
rect 582377 62781 582389 62784
rect 582423 62781 582435 62815
rect 582377 62775 582435 62781
rect 33042 62704 33048 62756
rect 33100 62744 33106 62756
rect 80330 62744 80336 62756
rect 33100 62716 80336 62744
rect 33100 62704 33106 62716
rect 80330 62704 80336 62716
rect 80388 62704 80394 62756
rect 80698 62704 80704 62756
rect 80756 62744 80762 62756
rect 90910 62744 90916 62756
rect 80756 62716 90916 62744
rect 80756 62704 80762 62716
rect 90910 62704 90916 62716
rect 90968 62704 90974 62756
rect 91738 62704 91744 62756
rect 91796 62744 91802 62756
rect 108298 62744 108304 62756
rect 91796 62716 108304 62744
rect 91796 62704 91802 62716
rect 108298 62704 108304 62716
rect 108356 62704 108362 62756
rect 117222 62704 117228 62756
rect 117280 62744 117286 62756
rect 148870 62744 148876 62756
rect 117280 62716 148876 62744
rect 117280 62704 117286 62716
rect 148870 62704 148876 62716
rect 148928 62704 148934 62756
rect 162762 62704 162768 62756
rect 162820 62744 162826 62756
rect 186590 62744 186596 62756
rect 162820 62716 186596 62744
rect 162820 62704 162826 62716
rect 186590 62704 186596 62716
rect 186648 62704 186654 62756
rect 188982 62704 188988 62756
rect 189040 62744 189046 62756
rect 207842 62744 207848 62756
rect 189040 62716 207848 62744
rect 189040 62704 189046 62716
rect 207842 62704 207848 62716
rect 207900 62704 207906 62756
rect 208302 62704 208308 62756
rect 208360 62744 208366 62756
rect 223298 62744 223304 62756
rect 208360 62716 223304 62744
rect 208360 62704 208366 62716
rect 223298 62704 223304 62716
rect 223356 62704 223362 62756
rect 235810 62704 235816 62756
rect 235868 62744 235874 62756
rect 245470 62744 245476 62756
rect 235868 62716 245476 62744
rect 235868 62704 235874 62716
rect 245470 62704 245476 62716
rect 245528 62704 245534 62756
rect 302510 62704 302516 62756
rect 302568 62744 302574 62756
rect 303338 62744 303344 62756
rect 302568 62716 303344 62744
rect 302568 62704 302574 62716
rect 303338 62704 303344 62716
rect 303396 62704 303402 62756
rect 325694 62704 325700 62756
rect 325752 62744 325758 62756
rect 331858 62744 331864 62756
rect 325752 62716 331864 62744
rect 325752 62704 325758 62716
rect 331858 62704 331864 62716
rect 331916 62704 331922 62756
rect 486050 62704 486056 62756
rect 486108 62744 486114 62756
rect 525058 62744 525064 62756
rect 486108 62716 525064 62744
rect 486108 62704 486114 62716
rect 525058 62704 525064 62716
rect 525116 62704 525122 62756
rect 528554 62704 528560 62756
rect 528612 62744 528618 62756
rect 545758 62744 545764 62756
rect 528612 62716 545764 62744
rect 528612 62704 528618 62716
rect 545758 62704 545764 62716
rect 545816 62704 545822 62756
rect 39942 62636 39948 62688
rect 40000 62676 40006 62688
rect 86126 62676 86132 62688
rect 40000 62648 86132 62676
rect 40000 62636 40006 62648
rect 86126 62636 86132 62648
rect 86184 62636 86190 62688
rect 122742 62636 122748 62688
rect 122800 62676 122806 62688
rect 153746 62676 153752 62688
rect 122800 62648 153752 62676
rect 122800 62636 122806 62648
rect 153746 62636 153752 62648
rect 153804 62636 153810 62688
rect 158622 62636 158628 62688
rect 158680 62676 158686 62688
rect 182726 62676 182732 62688
rect 158680 62648 182732 62676
rect 158680 62636 158686 62648
rect 182726 62636 182732 62648
rect 182784 62636 182790 62688
rect 190362 62636 190368 62688
rect 190420 62676 190426 62688
rect 208762 62676 208768 62688
rect 190420 62648 208768 62676
rect 190420 62636 190426 62648
rect 208762 62636 208768 62648
rect 208820 62636 208826 62688
rect 217962 62636 217968 62688
rect 218020 62676 218026 62688
rect 231026 62676 231032 62688
rect 218020 62648 231032 62676
rect 218020 62636 218026 62648
rect 231026 62636 231032 62648
rect 231084 62636 231090 62688
rect 313090 62636 313096 62688
rect 313148 62676 313154 62688
rect 313918 62676 313924 62688
rect 313148 62648 313924 62676
rect 313148 62636 313154 62648
rect 313918 62636 313924 62648
rect 313976 62636 313982 62688
rect 351730 62636 351736 62688
rect 351788 62676 351794 62688
rect 352558 62676 352564 62688
rect 351788 62648 352564 62676
rect 351788 62636 351794 62648
rect 352558 62636 352564 62648
rect 352616 62636 352622 62688
rect 487982 62636 487988 62688
rect 488040 62676 488046 62688
rect 526438 62676 526444 62688
rect 488040 62648 526444 62676
rect 488040 62636 488046 62648
rect 526438 62636 526444 62648
rect 526496 62636 526502 62688
rect 34422 62568 34428 62620
rect 34480 62608 34486 62620
rect 81250 62608 81256 62620
rect 34480 62580 81256 62608
rect 34480 62568 34486 62580
rect 81250 62568 81256 62580
rect 81308 62568 81314 62620
rect 97258 62568 97264 62620
rect 97316 62608 97322 62620
rect 106366 62608 106372 62620
rect 97316 62580 106372 62608
rect 97316 62568 97322 62580
rect 106366 62568 106372 62580
rect 106424 62568 106430 62620
rect 107010 62568 107016 62620
rect 107068 62608 107074 62620
rect 122834 62608 122840 62620
rect 107068 62580 122840 62608
rect 107068 62568 107074 62580
rect 122834 62568 122840 62580
rect 122892 62568 122898 62620
rect 125502 62568 125508 62620
rect 125560 62608 125566 62620
rect 155678 62608 155684 62620
rect 125560 62580 155684 62608
rect 125560 62568 125566 62580
rect 155678 62568 155684 62580
rect 155736 62568 155742 62620
rect 160002 62568 160008 62620
rect 160060 62608 160066 62620
rect 183646 62608 183652 62620
rect 160060 62580 183652 62608
rect 160060 62568 160066 62580
rect 183646 62568 183652 62580
rect 183704 62568 183710 62620
rect 184842 62568 184848 62620
rect 184900 62608 184906 62620
rect 203978 62608 203984 62620
rect 184900 62580 203984 62608
rect 184900 62568 184906 62580
rect 203978 62568 203984 62580
rect 204036 62568 204042 62620
rect 219342 62568 219348 62620
rect 219400 62608 219406 62620
rect 232958 62608 232964 62620
rect 219400 62580 232964 62608
rect 219400 62568 219406 62580
rect 232958 62568 232964 62580
rect 233016 62568 233022 62620
rect 452194 62568 452200 62620
rect 452252 62608 452258 62620
rect 453298 62608 453304 62620
rect 452252 62580 453304 62608
rect 452252 62568 452258 62580
rect 453298 62568 453304 62580
rect 453356 62568 453362 62620
rect 477310 62568 477316 62620
rect 477368 62608 477374 62620
rect 515490 62608 515496 62620
rect 477368 62580 515496 62608
rect 477368 62568 477374 62580
rect 515490 62568 515496 62580
rect 515548 62568 515554 62620
rect 515950 62568 515956 62620
rect 516008 62608 516014 62620
rect 517514 62608 517520 62620
rect 516008 62580 517520 62608
rect 516008 62568 516014 62580
rect 517514 62568 517520 62580
rect 517572 62568 517578 62620
rect 523678 62568 523684 62620
rect 523736 62608 523742 62620
rect 551278 62608 551284 62620
rect 523736 62580 551284 62608
rect 523736 62568 523742 62580
rect 551278 62568 551284 62580
rect 551336 62568 551342 62620
rect 41322 62500 41328 62552
rect 41380 62540 41386 62552
rect 87046 62540 87052 62552
rect 41380 62512 87052 62540
rect 41380 62500 41386 62512
rect 87046 62500 87052 62512
rect 87104 62500 87110 62552
rect 95878 62500 95884 62552
rect 95936 62540 95942 62552
rect 111242 62540 111248 62552
rect 95936 62512 111248 62540
rect 95936 62500 95942 62512
rect 111242 62500 111248 62512
rect 111300 62500 111306 62552
rect 116578 62500 116584 62552
rect 116636 62540 116642 62552
rect 143074 62540 143080 62552
rect 116636 62512 143080 62540
rect 116636 62500 116642 62512
rect 143074 62500 143080 62512
rect 143132 62500 143138 62552
rect 146938 62500 146944 62552
rect 146996 62540 147002 62552
rect 158530 62540 158536 62552
rect 146996 62512 158536 62540
rect 146996 62500 147002 62512
rect 158530 62500 158536 62512
rect 158588 62500 158594 62552
rect 164142 62500 164148 62552
rect 164200 62540 164206 62552
rect 187510 62540 187516 62552
rect 164200 62512 187516 62540
rect 164200 62500 164206 62512
rect 187510 62500 187516 62512
rect 187568 62500 187574 62552
rect 187602 62500 187608 62552
rect 187660 62540 187666 62552
rect 206830 62540 206836 62552
rect 187660 62512 206836 62540
rect 187660 62500 187666 62512
rect 206830 62500 206836 62512
rect 206888 62500 206894 62552
rect 216582 62500 216588 62552
rect 216640 62540 216646 62552
rect 230014 62540 230020 62552
rect 216640 62512 230020 62540
rect 216640 62500 216646 62512
rect 230014 62500 230020 62512
rect 230072 62500 230078 62552
rect 478322 62500 478328 62552
rect 478380 62540 478386 62552
rect 479518 62540 479524 62552
rect 478380 62512 479524 62540
rect 478380 62500 478386 62512
rect 479518 62500 479524 62512
rect 479576 62500 479582 62552
rect 513926 62540 513932 62552
rect 480226 62512 513932 62540
rect 50982 62432 50988 62484
rect 51040 62472 51046 62484
rect 94774 62472 94780 62484
rect 51040 62444 94780 62472
rect 51040 62432 51046 62444
rect 94774 62432 94780 62444
rect 94832 62432 94838 62484
rect 100110 62432 100116 62484
rect 100168 62472 100174 62484
rect 109310 62472 109316 62484
rect 100168 62444 109316 62472
rect 100168 62432 100174 62444
rect 109310 62432 109316 62444
rect 109368 62432 109374 62484
rect 112438 62432 112444 62484
rect 112496 62472 112502 62484
rect 128630 62472 128636 62484
rect 112496 62444 128636 62472
rect 112496 62432 112502 62444
rect 128630 62432 128636 62444
rect 128688 62432 128694 62484
rect 137278 62432 137284 62484
rect 137336 62472 137342 62484
rect 149882 62472 149888 62484
rect 137336 62444 149888 62472
rect 137336 62432 137342 62444
rect 149882 62432 149888 62444
rect 149940 62432 149946 62484
rect 161382 62432 161388 62484
rect 161440 62472 161446 62484
rect 184658 62472 184664 62484
rect 161440 62444 184664 62472
rect 161440 62432 161446 62444
rect 184658 62432 184664 62444
rect 184716 62432 184722 62484
rect 195882 62432 195888 62484
rect 195940 62472 195946 62484
rect 213638 62472 213644 62484
rect 195940 62444 213644 62472
rect 195940 62432 195946 62444
rect 213638 62432 213644 62444
rect 213696 62432 213702 62484
rect 321830 62432 321836 62484
rect 321888 62472 321894 62484
rect 322842 62472 322848 62484
rect 321888 62444 322848 62472
rect 321888 62432 321894 62444
rect 322842 62432 322848 62444
rect 322900 62432 322906 62484
rect 333422 62432 333428 62484
rect 333480 62472 333486 62484
rect 334618 62472 334624 62484
rect 333480 62444 334624 62472
rect 333480 62432 333486 62444
rect 334618 62432 334624 62444
rect 334676 62432 334682 62484
rect 391382 62432 391388 62484
rect 391440 62472 391446 62484
rect 392578 62472 392584 62484
rect 391440 62444 392584 62472
rect 391440 62432 391446 62444
rect 392578 62432 392584 62444
rect 392636 62432 392642 62484
rect 476390 62432 476396 62484
rect 476448 62472 476454 62484
rect 480226 62472 480254 62512
rect 513926 62500 513932 62512
rect 513984 62500 513990 62552
rect 519814 62500 519820 62552
rect 519872 62540 519878 62552
rect 534718 62540 534724 62552
rect 519872 62512 534724 62540
rect 519872 62500 519878 62512
rect 534718 62500 534724 62512
rect 534776 62500 534782 62552
rect 476448 62444 480254 62472
rect 476448 62432 476454 62444
rect 505370 62432 505376 62484
rect 505428 62472 505434 62484
rect 540330 62472 540336 62484
rect 505428 62444 540336 62472
rect 505428 62432 505434 62444
rect 540330 62432 540336 62444
rect 540388 62432 540394 62484
rect 43438 62364 43444 62416
rect 43496 62404 43502 62416
rect 79318 62404 79324 62416
rect 43496 62376 79324 62404
rect 43496 62364 43502 62376
rect 79318 62364 79324 62376
rect 79376 62364 79382 62416
rect 113818 62364 113824 62416
rect 113876 62404 113882 62416
rect 126698 62404 126704 62416
rect 113876 62376 126704 62404
rect 113876 62364 113882 62376
rect 126698 62364 126704 62376
rect 126756 62364 126762 62416
rect 135898 62364 135904 62416
rect 135956 62404 135962 62416
rect 146846 62404 146852 62416
rect 135956 62376 146852 62404
rect 135956 62364 135962 62376
rect 146846 62364 146852 62376
rect 146904 62364 146910 62416
rect 156598 62364 156604 62416
rect 156656 62404 156662 62416
rect 164326 62404 164332 62416
rect 156656 62376 164332 62404
rect 156656 62364 156662 62376
rect 164326 62364 164332 62376
rect 164384 62364 164390 62416
rect 166902 62364 166908 62416
rect 166960 62404 166966 62416
rect 189442 62404 189448 62416
rect 166960 62376 189448 62404
rect 166960 62364 166966 62376
rect 189442 62364 189448 62376
rect 189500 62364 189506 62416
rect 193122 62364 193128 62416
rect 193180 62404 193186 62416
rect 210694 62404 210700 62416
rect 193180 62376 210700 62404
rect 193180 62364 193186 62376
rect 210694 62364 210700 62376
rect 210752 62364 210758 62416
rect 260742 62364 260748 62416
rect 260800 62404 260806 62416
rect 266722 62404 266728 62416
rect 260800 62376 266728 62404
rect 260800 62364 260806 62376
rect 266722 62364 266728 62376
rect 266780 62364 266786 62416
rect 308306 62364 308312 62416
rect 308364 62404 308370 62416
rect 309778 62404 309784 62416
rect 308364 62376 309784 62404
rect 308364 62364 308370 62376
rect 309778 62364 309784 62376
rect 309836 62364 309842 62416
rect 341150 62364 341156 62416
rect 341208 62404 341214 62416
rect 342162 62404 342168 62416
rect 341208 62376 342168 62404
rect 341208 62364 341214 62376
rect 342162 62364 342168 62376
rect 342220 62364 342226 62416
rect 360470 62364 360476 62416
rect 360528 62404 360534 62416
rect 361482 62404 361488 62416
rect 360528 62376 361488 62404
rect 360528 62364 360534 62376
rect 361482 62364 361488 62376
rect 361540 62364 361546 62416
rect 399110 62364 399116 62416
rect 399168 62404 399174 62416
rect 400122 62404 400128 62416
rect 399168 62376 400128 62404
rect 399168 62364 399174 62376
rect 400122 62364 400128 62376
rect 400180 62364 400186 62416
rect 418430 62364 418436 62416
rect 418488 62404 418494 62416
rect 419442 62404 419448 62416
rect 418488 62376 419448 62404
rect 418488 62364 418494 62376
rect 419442 62364 419448 62376
rect 419500 62364 419506 62416
rect 420362 62364 420368 62416
rect 420420 62404 420426 62416
rect 421558 62404 421564 62416
rect 420420 62376 421564 62404
rect 420420 62364 420426 62376
rect 421558 62364 421564 62376
rect 421616 62364 421622 62416
rect 441614 62364 441620 62416
rect 441672 62404 441678 62416
rect 442902 62404 442908 62416
rect 441672 62376 442908 62404
rect 441672 62364 441678 62376
rect 442902 62364 442908 62376
rect 442960 62364 442966 62416
rect 483106 62364 483112 62416
rect 483164 62404 483170 62416
rect 515398 62404 515404 62416
rect 483164 62376 515404 62404
rect 483164 62364 483170 62376
rect 515398 62364 515404 62376
rect 515456 62364 515462 62416
rect 525610 62364 525616 62416
rect 525668 62404 525674 62416
rect 540238 62404 540244 62416
rect 525668 62376 540244 62404
rect 525668 62364 525674 62376
rect 540238 62364 540244 62376
rect 540296 62364 540302 62416
rect 53098 62296 53104 62348
rect 53156 62336 53162 62348
rect 93854 62336 93860 62348
rect 53156 62308 93860 62336
rect 53156 62296 53162 62308
rect 93854 62296 93860 62308
rect 93912 62296 93918 62348
rect 108298 62296 108304 62348
rect 108356 62336 108362 62348
rect 117958 62336 117964 62348
rect 108356 62308 117964 62336
rect 108356 62296 108362 62308
rect 117958 62296 117964 62308
rect 118016 62296 118022 62348
rect 123478 62296 123484 62348
rect 123536 62336 123542 62348
rect 135346 62336 135352 62348
rect 123536 62308 135352 62336
rect 123536 62296 123542 62308
rect 135346 62296 135352 62308
rect 135404 62296 135410 62348
rect 160738 62296 160744 62348
rect 160796 62336 160802 62348
rect 173066 62336 173072 62348
rect 160796 62308 173072 62336
rect 160796 62296 160802 62308
rect 173066 62296 173072 62308
rect 173124 62296 173130 62348
rect 173802 62296 173808 62348
rect 173860 62336 173866 62348
rect 195238 62336 195244 62348
rect 173860 62308 195244 62336
rect 173860 62296 173866 62308
rect 195238 62296 195244 62308
rect 195296 62296 195302 62348
rect 200022 62296 200028 62348
rect 200080 62336 200086 62348
rect 216490 62336 216496 62348
rect 200080 62308 216496 62336
rect 200080 62296 200086 62308
rect 216490 62296 216496 62308
rect 216548 62296 216554 62348
rect 259362 62296 259368 62348
rect 259420 62336 259426 62348
rect 264790 62336 264796 62348
rect 259420 62308 264796 62336
rect 259420 62296 259426 62308
rect 264790 62296 264796 62308
rect 264848 62296 264854 62348
rect 269022 62296 269028 62348
rect 269080 62336 269086 62348
rect 273530 62336 273536 62348
rect 269080 62308 273536 62336
rect 269080 62296 269086 62308
rect 273530 62296 273536 62308
rect 273588 62296 273594 62348
rect 316034 62296 316040 62348
rect 316092 62336 316098 62348
rect 317322 62336 317328 62348
rect 316092 62308 317328 62336
rect 316092 62296 316098 62308
rect 317322 62296 317328 62308
rect 317380 62296 317386 62348
rect 335354 62296 335360 62348
rect 335412 62336 335418 62348
rect 336642 62336 336648 62348
rect 335412 62308 336648 62336
rect 335412 62296 335418 62308
rect 336642 62296 336648 62308
rect 336700 62296 336706 62348
rect 338206 62296 338212 62348
rect 338264 62336 338270 62348
rect 339402 62336 339408 62348
rect 338264 62308 339408 62336
rect 338264 62296 338270 62308
rect 339402 62296 339408 62308
rect 339460 62296 339466 62348
rect 357526 62296 357532 62348
rect 357584 62336 357590 62348
rect 358722 62336 358728 62348
rect 357584 62308 358728 62336
rect 357584 62296 357590 62308
rect 358722 62296 358728 62308
rect 358780 62296 358786 62348
rect 373994 62296 374000 62348
rect 374052 62336 374058 62348
rect 375282 62336 375288 62348
rect 374052 62308 375288 62336
rect 374052 62296 374058 62308
rect 375282 62296 375288 62308
rect 375340 62296 375346 62348
rect 376846 62296 376852 62348
rect 376904 62336 376910 62348
rect 378042 62336 378048 62348
rect 376904 62308 378048 62336
rect 376904 62296 376910 62308
rect 378042 62296 378048 62308
rect 378100 62296 378106 62348
rect 379790 62296 379796 62348
rect 379848 62336 379854 62348
rect 381538 62336 381544 62348
rect 379848 62308 381544 62336
rect 379848 62296 379854 62308
rect 381538 62296 381544 62308
rect 381596 62296 381602 62348
rect 393314 62296 393320 62348
rect 393372 62336 393378 62348
rect 394602 62336 394608 62348
rect 393372 62308 394608 62336
rect 393372 62296 393378 62308
rect 394602 62296 394608 62308
rect 394660 62296 394666 62348
rect 396166 62296 396172 62348
rect 396224 62336 396230 62348
rect 397362 62336 397368 62348
rect 396224 62308 397368 62336
rect 396224 62296 396230 62308
rect 397362 62296 397368 62308
rect 397420 62296 397426 62348
rect 524690 62296 524696 62348
rect 524748 62336 524754 62348
rect 531958 62336 531964 62348
rect 524748 62308 531964 62336
rect 524748 62296 524754 62308
rect 531958 62296 531964 62308
rect 532016 62296 532022 62348
rect 15102 62228 15108 62280
rect 15160 62268 15166 62280
rect 65794 62268 65800 62280
rect 15160 62240 65800 62268
rect 15160 62228 15166 62240
rect 65794 62228 65800 62240
rect 65852 62228 65858 62280
rect 66898 62228 66904 62280
rect 66956 62268 66962 62280
rect 96706 62268 96712 62280
rect 66956 62240 96712 62268
rect 66956 62228 66962 62240
rect 96706 62228 96712 62240
rect 96764 62228 96770 62280
rect 98638 62228 98644 62280
rect 98696 62268 98702 62280
rect 114094 62268 114100 62280
rect 98696 62240 114100 62268
rect 98696 62228 98702 62240
rect 114094 62228 114100 62240
rect 114152 62228 114158 62280
rect 120718 62228 120724 62280
rect 120776 62268 120782 62280
rect 132494 62268 132500 62280
rect 120776 62240 132500 62268
rect 120776 62228 120782 62240
rect 132494 62228 132500 62240
rect 132552 62228 132558 62280
rect 176562 62228 176568 62280
rect 176620 62268 176626 62280
rect 197170 62268 197176 62280
rect 176620 62240 197176 62268
rect 176620 62228 176626 62240
rect 197170 62228 197176 62240
rect 197228 62228 197234 62280
rect 201402 62228 201408 62280
rect 201460 62268 201466 62280
rect 217502 62268 217508 62280
rect 201460 62240 217508 62268
rect 201460 62228 201466 62240
rect 217502 62228 217508 62240
rect 217560 62228 217566 62280
rect 249702 62228 249708 62280
rect 249760 62268 249766 62280
rect 257062 62268 257068 62280
rect 249760 62240 257068 62268
rect 249760 62228 249766 62240
rect 257062 62228 257068 62240
rect 257120 62228 257126 62280
rect 263502 62228 263508 62280
rect 263560 62268 263566 62280
rect 268654 62268 268660 62280
rect 263560 62240 268660 62268
rect 263560 62228 263566 62240
rect 268654 62228 268660 62240
rect 268712 62228 268718 62280
rect 270402 62228 270408 62280
rect 270460 62268 270466 62280
rect 274450 62268 274456 62280
rect 270460 62240 274456 62268
rect 270460 62228 270466 62240
rect 274450 62228 274456 62240
rect 274508 62228 274514 62280
rect 274542 62228 274548 62280
rect 274600 62268 274606 62280
rect 277394 62268 277400 62280
rect 274600 62240 277400 62268
rect 274600 62228 274606 62240
rect 277394 62228 277400 62240
rect 277452 62228 277458 62280
rect 319898 62228 319904 62280
rect 319956 62268 319962 62280
rect 320910 62268 320916 62280
rect 319956 62240 320916 62268
rect 319956 62228 319962 62240
rect 320910 62228 320916 62240
rect 320968 62228 320974 62280
rect 408770 62228 408776 62280
rect 408828 62268 408834 62280
rect 410518 62268 410524 62280
rect 408828 62240 410524 62268
rect 408828 62228 408834 62240
rect 410518 62228 410524 62240
rect 410576 62228 410582 62280
rect 450262 62228 450268 62280
rect 450320 62268 450326 62280
rect 451182 62268 451188 62280
rect 450320 62240 451188 62268
rect 450320 62228 450326 62240
rect 451182 62228 451188 62240
rect 451240 62228 451246 62280
rect 481174 62228 481180 62280
rect 481232 62268 481238 62280
rect 485130 62268 485136 62280
rect 481232 62240 485136 62268
rect 481232 62228 481238 62240
rect 485130 62228 485136 62240
rect 485188 62228 485194 62280
rect 55858 62160 55864 62212
rect 55916 62200 55922 62212
rect 84194 62200 84200 62212
rect 55916 62172 84200 62200
rect 55916 62160 55922 62172
rect 84194 62160 84200 62172
rect 84252 62160 84258 62212
rect 106918 62160 106924 62212
rect 106976 62200 106982 62212
rect 115106 62200 115112 62212
rect 106976 62172 115112 62200
rect 106976 62160 106982 62172
rect 115106 62160 115112 62172
rect 115164 62160 115170 62212
rect 133138 62160 133144 62212
rect 133196 62200 133202 62212
rect 141142 62200 141148 62212
rect 133196 62172 141148 62200
rect 133196 62160 133202 62172
rect 141142 62160 141148 62172
rect 141200 62160 141206 62212
rect 188338 62160 188344 62212
rect 188396 62200 188402 62212
rect 204898 62200 204904 62212
rect 188396 62172 204904 62200
rect 188396 62160 188402 62172
rect 204898 62160 204904 62172
rect 204956 62160 204962 62212
rect 252370 62160 252376 62212
rect 252428 62200 252434 62212
rect 260006 62200 260012 62212
rect 252428 62172 260012 62200
rect 252428 62160 252434 62172
rect 260006 62160 260012 62172
rect 260064 62160 260070 62212
rect 264882 62160 264888 62212
rect 264940 62200 264946 62212
rect 269666 62200 269672 62212
rect 264940 62172 269672 62200
rect 264940 62160 264946 62172
rect 269666 62160 269672 62172
rect 269724 62160 269730 62212
rect 271782 62160 271788 62212
rect 271840 62200 271846 62212
rect 275462 62200 275468 62212
rect 271840 62172 275468 62200
rect 271840 62160 271846 62172
rect 275462 62160 275468 62172
rect 275520 62160 275526 62212
rect 275922 62160 275928 62212
rect 275980 62200 275986 62212
rect 278314 62200 278320 62212
rect 275980 62172 278320 62200
rect 275980 62160 275986 62172
rect 278314 62160 278320 62172
rect 278372 62160 278378 62212
rect 278682 62160 278688 62212
rect 278740 62200 278746 62212
rect 281258 62200 281264 62212
rect 278740 62172 281264 62200
rect 278740 62160 278746 62172
rect 281258 62160 281264 62172
rect 281316 62160 281322 62212
rect 281442 62160 281448 62212
rect 281500 62200 281506 62212
rect 283190 62200 283196 62212
rect 281500 62172 283196 62200
rect 281500 62160 281506 62172
rect 283190 62160 283196 62172
rect 283248 62160 283254 62212
rect 315022 62160 315028 62212
rect 315080 62200 315086 62212
rect 318058 62200 318064 62212
rect 315080 62172 318064 62200
rect 315080 62160 315086 62172
rect 318058 62160 318064 62172
rect 318116 62160 318122 62212
rect 433886 62160 433892 62212
rect 433944 62200 433950 62212
rect 439498 62200 439504 62212
rect 433944 62172 439504 62200
rect 433944 62160 433950 62172
rect 439498 62160 439504 62172
rect 439556 62160 439562 62212
rect 469582 62160 469588 62212
rect 469640 62200 469646 62212
rect 472618 62200 472624 62212
rect 469640 62172 472624 62200
rect 469640 62160 469646 62172
rect 472618 62160 472624 62172
rect 472676 62160 472682 62212
rect 473446 62160 473452 62212
rect 473504 62200 473510 62212
rect 476758 62200 476764 62212
rect 473504 62172 476764 62200
rect 473504 62160 473510 62172
rect 476758 62160 476764 62172
rect 476816 62160 476822 62212
rect 480254 62160 480260 62212
rect 480312 62200 480318 62212
rect 483658 62200 483664 62212
rect 480312 62172 483664 62200
rect 480312 62160 480318 62172
rect 483658 62160 483664 62172
rect 483716 62160 483722 62212
rect 510154 62160 510160 62212
rect 510212 62200 510218 62212
rect 511258 62200 511264 62212
rect 510212 62172 511264 62200
rect 510212 62160 510218 62172
rect 511258 62160 511264 62172
rect 511316 62160 511322 62212
rect 59998 62092 60004 62144
rect 60056 62132 60062 62144
rect 61010 62132 61016 62144
rect 60056 62104 61016 62132
rect 60056 62092 60062 62104
rect 61010 62092 61016 62104
rect 61068 62092 61074 62144
rect 61378 62092 61384 62144
rect 61436 62132 61442 62144
rect 75089 62135 75147 62141
rect 75089 62132 75101 62135
rect 61436 62104 75101 62132
rect 61436 62092 61442 62104
rect 75089 62101 75101 62104
rect 75135 62101 75147 62135
rect 75089 62095 75147 62101
rect 75178 62092 75184 62144
rect 75236 62132 75242 62144
rect 82262 62132 82268 62144
rect 75236 62104 82268 62132
rect 75236 62092 75242 62104
rect 82262 62092 82268 62104
rect 82320 62092 82326 62144
rect 88978 62092 88984 62144
rect 89036 62132 89042 62144
rect 91922 62132 91928 62144
rect 89036 62104 91928 62132
rect 89036 62092 89042 62104
rect 91922 62092 91928 62104
rect 91980 62092 91986 62144
rect 100018 62092 100024 62144
rect 100076 62132 100082 62144
rect 103514 62132 103520 62144
rect 100076 62104 103520 62132
rect 100076 62092 100082 62104
rect 103514 62092 103520 62104
rect 103572 62092 103578 62144
rect 113910 62092 113916 62144
rect 113968 62132 113974 62144
rect 120902 62132 120908 62144
rect 113968 62104 120908 62132
rect 113968 62092 113974 62104
rect 120902 62092 120908 62104
rect 120960 62092 120966 62144
rect 134610 62092 134616 62144
rect 134668 62132 134674 62144
rect 136358 62132 136364 62144
rect 134668 62104 136364 62132
rect 134668 62092 134674 62104
rect 136358 62092 136364 62104
rect 136416 62092 136422 62144
rect 137370 62092 137376 62144
rect 137428 62132 137434 62144
rect 139210 62132 139216 62144
rect 137428 62104 139216 62132
rect 137428 62092 137434 62104
rect 139210 62092 139216 62104
rect 139268 62092 139274 62144
rect 202782 62092 202788 62144
rect 202840 62132 202846 62144
rect 218422 62132 218428 62144
rect 202840 62104 218428 62132
rect 202840 62092 202846 62104
rect 218422 62092 218428 62104
rect 218480 62092 218486 62144
rect 252462 62092 252468 62144
rect 252520 62132 252526 62144
rect 258994 62132 259000 62144
rect 252520 62104 259000 62132
rect 252520 62092 252526 62104
rect 258994 62092 259000 62104
rect 259052 62092 259058 62144
rect 260650 62092 260656 62144
rect 260708 62132 260714 62144
rect 265802 62132 265808 62144
rect 260708 62104 265808 62132
rect 260708 62092 260714 62104
rect 265802 62092 265808 62104
rect 265860 62092 265866 62144
rect 267090 62092 267096 62144
rect 267148 62132 267154 62144
rect 267734 62132 267740 62144
rect 267148 62104 267740 62132
rect 267148 62092 267154 62104
rect 267734 62092 267740 62104
rect 267792 62092 267798 62144
rect 269758 62092 269764 62144
rect 269816 62132 269822 62144
rect 272518 62132 272524 62144
rect 269816 62104 272524 62132
rect 269816 62092 269822 62104
rect 272518 62092 272524 62104
rect 272576 62092 272582 62144
rect 277302 62092 277308 62144
rect 277360 62132 277366 62144
rect 279326 62132 279332 62144
rect 277360 62104 279332 62132
rect 277360 62092 277366 62104
rect 279326 62092 279332 62104
rect 279384 62092 279390 62144
rect 280798 62092 280804 62144
rect 280856 62132 280862 62144
rect 282178 62132 282184 62144
rect 280856 62104 282184 62132
rect 280856 62092 280862 62104
rect 282178 62092 282184 62104
rect 282236 62092 282242 62144
rect 282822 62092 282828 62144
rect 282880 62132 282886 62144
rect 284110 62132 284116 62144
rect 282880 62104 284116 62132
rect 282880 62092 282886 62104
rect 284110 62092 284116 62104
rect 284168 62092 284174 62144
rect 285582 62092 285588 62144
rect 285640 62132 285646 62144
rect 287054 62132 287060 62144
rect 285640 62104 287060 62132
rect 285640 62092 285646 62104
rect 287054 62092 287060 62104
rect 287112 62092 287118 62144
rect 288342 62092 288348 62144
rect 288400 62132 288406 62144
rect 288986 62132 288992 62144
rect 288400 62104 288992 62132
rect 288400 62092 288406 62104
rect 288986 62092 288992 62104
rect 289044 62092 289050 62144
rect 289814 62092 289820 62144
rect 289872 62132 289878 62144
rect 290918 62132 290924 62144
rect 289872 62104 290924 62132
rect 289872 62092 289878 62104
rect 290918 62092 290924 62104
rect 290976 62092 290982 62144
rect 292574 62092 292580 62144
rect 292632 62132 292638 62144
rect 293770 62132 293776 62144
rect 292632 62104 293776 62132
rect 292632 62092 292638 62104
rect 293770 62092 293776 62104
rect 293828 62092 293834 62144
rect 297634 62092 297640 62144
rect 297692 62132 297698 62144
rect 298186 62132 298192 62144
rect 297692 62104 298192 62132
rect 297692 62092 297698 62104
rect 298186 62092 298192 62104
rect 298244 62092 298250 62144
rect 298646 62092 298652 62144
rect 298704 62132 298710 62144
rect 299382 62132 299388 62144
rect 298704 62104 299388 62132
rect 298704 62092 298710 62104
rect 299382 62092 299388 62104
rect 299440 62092 299446 62144
rect 301498 62092 301504 62144
rect 301556 62132 301562 62144
rect 302418 62132 302424 62144
rect 301556 62104 302424 62132
rect 301556 62092 301562 62104
rect 302418 62092 302424 62104
rect 302476 62092 302482 62144
rect 304442 62092 304448 62144
rect 304500 62132 304506 62144
rect 304902 62132 304908 62144
rect 304500 62104 304908 62132
rect 304500 62092 304506 62104
rect 304902 62092 304908 62104
rect 304960 62092 304966 62144
rect 305362 62092 305368 62144
rect 305420 62132 305426 62144
rect 306282 62132 306288 62144
rect 305420 62104 306288 62132
rect 305420 62092 305426 62104
rect 306282 62092 306288 62104
rect 306340 62092 306346 62144
rect 306374 62092 306380 62144
rect 306432 62132 306438 62144
rect 307662 62132 307668 62144
rect 306432 62104 307668 62132
rect 306432 62092 306438 62104
rect 307662 62092 307668 62104
rect 307720 62092 307726 62144
rect 309226 62092 309232 62144
rect 309284 62132 309290 62144
rect 310330 62132 310336 62144
rect 309284 62104 310336 62132
rect 309284 62092 309290 62104
rect 310330 62092 310336 62104
rect 310388 62092 310394 62144
rect 312170 62092 312176 62144
rect 312228 62132 312234 62144
rect 313182 62132 313188 62144
rect 312228 62104 313188 62132
rect 312228 62092 312234 62104
rect 313182 62092 313188 62104
rect 313240 62092 313246 62144
rect 314102 62092 314108 62144
rect 314160 62132 314166 62144
rect 314562 62132 314568 62144
rect 314160 62104 314568 62132
rect 314160 62092 314166 62104
rect 314562 62092 314568 62104
rect 314620 62092 314626 62144
rect 317966 62092 317972 62144
rect 318024 62132 318030 62144
rect 318702 62132 318708 62144
rect 318024 62104 318708 62132
rect 318024 62092 318030 62104
rect 318702 62092 318708 62104
rect 318760 62092 318766 62144
rect 320818 62092 320824 62144
rect 320876 62132 320882 62144
rect 321462 62132 321468 62144
rect 320876 62104 321468 62132
rect 320876 62092 320882 62104
rect 321462 62092 321468 62104
rect 321520 62092 321526 62144
rect 323762 62092 323768 62144
rect 323820 62132 323826 62144
rect 324222 62132 324228 62144
rect 323820 62104 324228 62132
rect 323820 62092 323826 62104
rect 324222 62092 324228 62104
rect 324280 62092 324286 62144
rect 324682 62092 324688 62144
rect 324740 62132 324746 62144
rect 325602 62132 325608 62144
rect 324740 62104 325608 62132
rect 324740 62092 324746 62104
rect 325602 62092 325608 62104
rect 325660 62092 325666 62144
rect 331490 62092 331496 62144
rect 331548 62132 331554 62144
rect 332318 62132 332324 62144
rect 331548 62104 332324 62132
rect 331548 62092 331554 62104
rect 332318 62092 332324 62104
rect 332376 62092 332382 62144
rect 337286 62092 337292 62144
rect 337344 62132 337350 62144
rect 340230 62132 340236 62144
rect 337344 62104 340236 62132
rect 337344 62092 337350 62104
rect 340230 62092 340236 62104
rect 340288 62092 340294 62144
rect 343082 62092 343088 62144
rect 343140 62132 343146 62144
rect 343542 62132 343548 62144
rect 343140 62104 343548 62132
rect 343140 62092 343146 62104
rect 343542 62092 343548 62104
rect 343600 62092 343606 62144
rect 344002 62092 344008 62144
rect 344060 62132 344066 62144
rect 344922 62132 344928 62144
rect 344060 62104 344928 62132
rect 344060 62092 344066 62104
rect 344922 62092 344928 62104
rect 344980 62092 344986 62144
rect 345014 62092 345020 62144
rect 345072 62132 345078 62144
rect 346210 62132 346216 62144
rect 345072 62104 346216 62132
rect 345072 62092 345078 62104
rect 346210 62092 346216 62104
rect 346268 62092 346274 62144
rect 347866 62092 347872 62144
rect 347924 62132 347930 62144
rect 349062 62132 349068 62144
rect 347924 62104 349068 62132
rect 347924 62092 347930 62104
rect 349062 62092 349068 62104
rect 349120 62092 349126 62144
rect 350810 62092 350816 62144
rect 350868 62132 350874 62144
rect 351822 62132 351828 62144
rect 350868 62104 351828 62132
rect 350868 62092 350874 62104
rect 351822 62092 351828 62104
rect 351880 62092 351886 62144
rect 352742 62092 352748 62144
rect 352800 62132 352806 62144
rect 353202 62132 353208 62144
rect 352800 62104 353208 62132
rect 352800 62092 352806 62104
rect 353202 62092 353208 62104
rect 353260 62092 353266 62144
rect 354674 62092 354680 62144
rect 354732 62132 354738 62144
rect 355870 62132 355876 62144
rect 354732 62104 355876 62132
rect 354732 62092 354738 62104
rect 355870 62092 355876 62104
rect 355928 62092 355934 62144
rect 356606 62092 356612 62144
rect 356664 62132 356670 62144
rect 357342 62132 357348 62144
rect 356664 62104 357348 62132
rect 356664 62092 356670 62104
rect 357342 62092 357348 62104
rect 357400 62092 357406 62144
rect 362402 62092 362408 62144
rect 362460 62132 362466 62144
rect 362862 62132 362868 62144
rect 362460 62104 362868 62132
rect 362460 62092 362466 62104
rect 362862 62092 362868 62104
rect 362920 62092 362926 62144
rect 363322 62092 363328 62144
rect 363380 62132 363386 62144
rect 364242 62132 364248 62144
rect 363380 62104 364248 62132
rect 363380 62092 363386 62104
rect 364242 62092 364248 62104
rect 364300 62092 364306 62144
rect 364334 62092 364340 62144
rect 364392 62132 364398 62144
rect 365622 62132 365628 62144
rect 364392 62104 365628 62132
rect 364392 62092 364398 62104
rect 365622 62092 365628 62104
rect 365680 62092 365686 62144
rect 370130 62092 370136 62144
rect 370188 62132 370194 62144
rect 371142 62132 371148 62144
rect 370188 62104 371148 62132
rect 370188 62092 370194 62104
rect 371142 62092 371148 62104
rect 371200 62092 371206 62144
rect 372062 62092 372068 62144
rect 372120 62132 372126 62144
rect 372522 62132 372528 62144
rect 372120 62104 372528 62132
rect 372120 62092 372126 62104
rect 372522 62092 372528 62104
rect 372580 62092 372586 62144
rect 375926 62092 375932 62144
rect 375984 62132 375990 62144
rect 376662 62132 376668 62144
rect 375984 62104 376668 62132
rect 375984 62092 375990 62104
rect 376662 62092 376668 62104
rect 376720 62092 376726 62144
rect 381722 62092 381728 62144
rect 381780 62132 381786 62144
rect 382182 62132 382188 62144
rect 381780 62104 382188 62132
rect 381780 62092 381786 62104
rect 382182 62092 382188 62104
rect 382240 62092 382246 62144
rect 382642 62092 382648 62144
rect 382700 62132 382706 62144
rect 383562 62132 383568 62144
rect 382700 62104 383568 62132
rect 382700 62092 382706 62104
rect 383562 62092 383568 62104
rect 383620 62092 383626 62144
rect 383654 62092 383660 62144
rect 383712 62132 383718 62144
rect 384850 62132 384856 62144
rect 383712 62104 384856 62132
rect 383712 62092 383718 62104
rect 384850 62092 384856 62104
rect 384908 62092 384914 62144
rect 389450 62092 389456 62144
rect 389508 62132 389514 62144
rect 390278 62132 390284 62144
rect 389508 62104 390284 62132
rect 389508 62092 389514 62104
rect 390278 62092 390284 62104
rect 390336 62092 390342 62144
rect 395246 62092 395252 62144
rect 395304 62132 395310 62144
rect 395982 62132 395988 62144
rect 395304 62104 395988 62132
rect 395304 62092 395310 62104
rect 395982 62092 395988 62104
rect 396040 62092 396046 62144
rect 401042 62092 401048 62144
rect 401100 62132 401106 62144
rect 401502 62132 401508 62144
rect 401100 62104 401508 62132
rect 401100 62092 401106 62104
rect 401502 62092 401508 62104
rect 401560 62092 401566 62144
rect 401962 62092 401968 62144
rect 402020 62132 402026 62144
rect 402882 62132 402888 62144
rect 402020 62104 402888 62132
rect 402020 62092 402026 62104
rect 402882 62092 402888 62104
rect 402940 62092 402946 62144
rect 402974 62092 402980 62144
rect 403032 62132 403038 62144
rect 404170 62132 404176 62144
rect 403032 62104 404176 62132
rect 403032 62092 403038 62104
rect 404170 62092 404176 62104
rect 404228 62092 404234 62144
rect 410702 62092 410708 62144
rect 410760 62132 410766 62144
rect 411162 62132 411168 62144
rect 410760 62104 411168 62132
rect 410760 62092 410766 62104
rect 411162 62092 411168 62104
rect 411220 62092 411226 62144
rect 412634 62092 412640 62144
rect 412692 62132 412698 62144
rect 413830 62132 413836 62144
rect 412692 62104 413836 62132
rect 412692 62092 412698 62104
rect 413830 62092 413836 62104
rect 413888 62092 413894 62144
rect 414566 62092 414572 62144
rect 414624 62132 414630 62144
rect 415302 62132 415308 62144
rect 414624 62104 415308 62132
rect 414624 62092 414630 62104
rect 415302 62092 415308 62104
rect 415360 62092 415366 62144
rect 415486 62092 415492 62144
rect 415544 62132 415550 62144
rect 416682 62132 416688 62144
rect 415544 62104 416688 62132
rect 415544 62092 415550 62104
rect 416682 62092 416688 62104
rect 416740 62092 416746 62144
rect 425146 62092 425152 62144
rect 425204 62132 425210 62144
rect 426342 62132 426348 62144
rect 425204 62104 426348 62132
rect 425204 62092 425210 62104
rect 426342 62092 426348 62104
rect 426400 62092 426406 62144
rect 428090 62092 428096 62144
rect 428148 62132 428154 62144
rect 429102 62132 429108 62144
rect 428148 62104 429108 62132
rect 428148 62092 428154 62104
rect 429102 62092 429108 62104
rect 429160 62092 429166 62144
rect 430022 62092 430028 62144
rect 430080 62132 430086 62144
rect 430482 62132 430488 62144
rect 430080 62104 430488 62132
rect 430080 62092 430086 62104
rect 430482 62092 430488 62104
rect 430540 62092 430546 62144
rect 430942 62092 430948 62144
rect 431000 62132 431006 62144
rect 431862 62132 431868 62144
rect 431000 62104 431868 62132
rect 431000 62092 431006 62104
rect 431862 62092 431868 62104
rect 431920 62092 431926 62144
rect 431954 62092 431960 62144
rect 432012 62132 432018 62144
rect 433150 62132 433156 62144
rect 432012 62104 433156 62132
rect 432012 62092 432018 62104
rect 433150 62092 433156 62104
rect 433208 62092 433214 62144
rect 436738 62092 436744 62144
rect 436796 62132 436802 62144
rect 437382 62132 437388 62144
rect 436796 62104 437388 62132
rect 436796 62092 436802 62104
rect 437382 62092 437388 62104
rect 437440 62092 437446 62144
rect 443546 62092 443552 62144
rect 443604 62132 443610 62144
rect 444282 62132 444288 62144
rect 443604 62104 444288 62132
rect 443604 62092 443610 62104
rect 444282 62092 444288 62104
rect 444340 62092 444346 62144
rect 446398 62092 446404 62144
rect 446456 62132 446462 62144
rect 447042 62132 447048 62144
rect 446456 62104 447048 62132
rect 446456 62092 446462 62104
rect 447042 62092 447048 62104
rect 447100 62092 447106 62144
rect 447410 62092 447416 62144
rect 447468 62132 447474 62144
rect 448238 62132 448244 62144
rect 447468 62104 448244 62132
rect 447468 62092 447474 62104
rect 448238 62092 448244 62104
rect 448296 62092 448302 62144
rect 449342 62092 449348 62144
rect 449400 62132 449406 62144
rect 449802 62132 449808 62144
rect 449400 62104 449808 62132
rect 449400 62092 449406 62104
rect 449802 62092 449808 62104
rect 449860 62092 449866 62144
rect 453206 62092 453212 62144
rect 453264 62132 453270 62144
rect 453942 62132 453948 62144
rect 453264 62104 453948 62132
rect 453264 62092 453270 62104
rect 453942 62092 453948 62104
rect 454000 62092 454006 62144
rect 456058 62092 456064 62144
rect 456116 62132 456122 62144
rect 456702 62132 456708 62144
rect 456116 62104 456708 62132
rect 456116 62092 456122 62104
rect 456702 62092 456708 62104
rect 456760 62092 456766 62144
rect 459002 62092 459008 62144
rect 459060 62132 459066 62144
rect 459462 62132 459468 62144
rect 459060 62104 459468 62132
rect 459060 62092 459066 62104
rect 459462 62092 459468 62104
rect 459520 62092 459526 62144
rect 459922 62092 459928 62144
rect 459980 62132 459986 62144
rect 460842 62132 460848 62144
rect 459980 62104 460848 62132
rect 459980 62092 459986 62104
rect 460842 62092 460848 62104
rect 460900 62092 460906 62144
rect 460934 62092 460940 62144
rect 460992 62132 460998 62144
rect 462130 62132 462136 62144
rect 460992 62104 462136 62132
rect 460992 62092 460998 62104
rect 462130 62092 462136 62104
rect 462188 62092 462194 62144
rect 465718 62092 465724 62144
rect 465776 62132 465782 62144
rect 466362 62132 466368 62144
rect 465776 62104 466368 62132
rect 465776 62092 465782 62104
rect 466362 62092 466368 62104
rect 466420 62092 466426 62144
rect 466730 62092 466736 62144
rect 466788 62132 466794 62144
rect 467742 62132 467748 62144
rect 466788 62104 467748 62132
rect 466788 62092 466794 62104
rect 467742 62092 467748 62104
rect 467800 62092 467806 62144
rect 472526 62092 472532 62144
rect 472584 62132 472590 62144
rect 473262 62132 473268 62144
rect 472584 62104 473268 62132
rect 472584 62092 472590 62104
rect 473262 62092 473268 62104
rect 473320 62092 473326 62144
rect 475378 62092 475384 62144
rect 475436 62132 475442 62144
rect 476022 62132 476028 62144
rect 475436 62104 476028 62132
rect 475436 62092 475442 62104
rect 476022 62092 476028 62104
rect 476080 62092 476086 62144
rect 479242 62092 479248 62144
rect 479300 62132 479306 62144
rect 480162 62132 480168 62144
rect 479300 62104 480168 62132
rect 479300 62092 479306 62104
rect 480162 62092 480168 62104
rect 480220 62092 480226 62144
rect 485038 62092 485044 62144
rect 485096 62132 485102 62144
rect 485682 62132 485688 62144
rect 485096 62104 485688 62132
rect 485096 62092 485102 62104
rect 485682 62092 485688 62104
rect 485740 62092 485746 62144
rect 488902 62092 488908 62144
rect 488960 62132 488966 62144
rect 489822 62132 489828 62144
rect 488960 62104 489828 62132
rect 488960 62092 488966 62104
rect 489822 62092 489828 62104
rect 489880 62092 489886 62144
rect 495710 62092 495716 62144
rect 495768 62132 495774 62144
rect 497550 62132 497556 62144
rect 495768 62104 497556 62132
rect 495768 62092 495774 62104
rect 497550 62092 497556 62104
rect 497608 62092 497614 62144
rect 498562 62092 498568 62144
rect 498620 62132 498626 62144
rect 500218 62132 500224 62144
rect 498620 62104 500224 62132
rect 498620 62092 498626 62104
rect 500218 62092 500224 62104
rect 500276 62092 500282 62144
rect 501506 62092 501512 62144
rect 501564 62132 501570 62144
rect 502242 62132 502248 62144
rect 501564 62104 502248 62132
rect 501564 62092 501570 62104
rect 502242 62092 502248 62104
rect 502300 62092 502306 62144
rect 502426 62092 502432 62144
rect 502484 62132 502490 62144
rect 503622 62132 503628 62144
rect 502484 62104 503628 62132
rect 502484 62092 502490 62104
rect 503622 62092 503628 62104
rect 503680 62092 503686 62144
rect 504358 62092 504364 62144
rect 504416 62132 504422 62144
rect 505002 62132 505008 62144
rect 504416 62104 505008 62132
rect 504416 62092 504422 62104
rect 505002 62092 505008 62104
rect 505060 62092 505066 62144
rect 507302 62092 507308 62144
rect 507360 62132 507366 62144
rect 507762 62132 507768 62144
rect 507360 62104 507768 62132
rect 507360 62092 507366 62104
rect 507762 62092 507768 62104
rect 507820 62092 507826 62144
rect 508222 62092 508228 62144
rect 508280 62132 508286 62144
rect 509142 62132 509148 62144
rect 508280 62104 509148 62132
rect 508280 62092 508286 62104
rect 509142 62092 509148 62104
rect 509200 62092 509206 62144
rect 511166 62092 511172 62144
rect 511224 62132 511230 62144
rect 511902 62132 511908 62144
rect 511224 62104 511908 62132
rect 511224 62092 511230 62104
rect 511902 62092 511908 62104
rect 511960 62092 511966 62144
rect 512086 62092 512092 62144
rect 512144 62132 512150 62144
rect 513190 62132 513196 62144
rect 512144 62104 513196 62132
rect 512144 62092 512150 62104
rect 513190 62092 513196 62104
rect 513248 62092 513254 62144
rect 514018 62092 514024 62144
rect 514076 62132 514082 62144
rect 514662 62132 514668 62144
rect 514076 62104 514668 62132
rect 514076 62092 514082 62104
rect 514662 62092 514668 62104
rect 514720 62092 514726 62144
rect 515030 62092 515036 62144
rect 515088 62132 515094 62144
rect 516042 62132 516048 62144
rect 515088 62104 516048 62132
rect 515088 62092 515094 62104
rect 516042 62092 516048 62104
rect 516100 62092 516106 62144
rect 516962 62092 516968 62144
rect 517020 62132 517026 62144
rect 517422 62132 517428 62144
rect 517020 62104 517428 62132
rect 517020 62092 517026 62104
rect 517422 62092 517428 62104
rect 517480 62092 517486 62144
rect 517882 62092 517888 62144
rect 517940 62132 517946 62144
rect 518802 62132 518808 62144
rect 517940 62104 518808 62132
rect 517940 62092 517946 62104
rect 518802 62092 518808 62104
rect 518860 62092 518866 62144
rect 518894 62092 518900 62144
rect 518952 62132 518958 62144
rect 520182 62132 520188 62144
rect 518952 62104 520188 62132
rect 518952 62092 518958 62104
rect 520182 62092 520188 62104
rect 520240 62092 520246 62144
rect 520826 62092 520832 62144
rect 520884 62132 520890 62144
rect 521562 62132 521568 62144
rect 520884 62104 521568 62132
rect 520884 62092 520890 62104
rect 521562 62092 521568 62104
rect 521620 62092 521626 62144
rect 526622 62092 526628 62144
rect 526680 62132 526686 62144
rect 527082 62132 527088 62144
rect 526680 62104 527088 62132
rect 526680 62092 526686 62104
rect 527082 62092 527088 62104
rect 527140 62092 527146 62144
rect 527542 62092 527548 62144
rect 527600 62132 527606 62144
rect 528462 62132 528468 62144
rect 527600 62104 528468 62132
rect 527600 62092 527606 62104
rect 528462 62092 528468 62104
rect 528520 62092 528526 62144
rect 36538 61956 36544 62008
rect 36596 61996 36602 62008
rect 55214 61996 55220 62008
rect 36596 61968 55220 61996
rect 36596 61956 36602 61968
rect 55214 61956 55220 61968
rect 55272 61956 55278 62008
rect 91002 61956 91008 62008
rect 91060 61996 91066 62008
rect 127618 61996 127624 62008
rect 91060 61968 127624 61996
rect 91060 61956 91066 61968
rect 127618 61956 127624 61968
rect 127676 61956 127682 62008
rect 151078 61956 151084 62008
rect 151136 61996 151142 62008
rect 162394 61996 162400 62008
rect 151136 61968 162400 61996
rect 151136 61956 151142 61968
rect 162394 61956 162400 61968
rect 162452 61956 162458 62008
rect 29730 61888 29736 61940
rect 29788 61928 29794 61940
rect 63862 61928 63868 61940
rect 29788 61900 63868 61928
rect 29788 61888 29794 61900
rect 63862 61888 63868 61900
rect 63920 61888 63926 61940
rect 84102 61888 84108 61940
rect 84160 61928 84166 61940
rect 121822 61928 121828 61940
rect 84160 61900 121828 61928
rect 84160 61888 84166 61900
rect 121822 61888 121828 61900
rect 121880 61888 121886 61940
rect 141418 61888 141424 61940
rect 141476 61928 141482 61940
rect 165338 61928 165344 61940
rect 141476 61900 165344 61928
rect 141476 61888 141482 61900
rect 165338 61888 165344 61900
rect 165396 61888 165402 61940
rect 35250 61820 35256 61872
rect 35308 61860 35314 61872
rect 75454 61860 75460 61872
rect 35308 61832 75460 61860
rect 35308 61820 35314 61832
rect 75454 61820 75460 61832
rect 75512 61820 75518 61872
rect 79962 61820 79968 61872
rect 80020 61860 80026 61872
rect 118970 61860 118976 61872
rect 80020 61832 118976 61860
rect 80020 61820 80026 61832
rect 118970 61820 118976 61832
rect 119028 61820 119034 61872
rect 151722 61820 151728 61872
rect 151780 61860 151786 61872
rect 176930 61860 176936 61872
rect 151780 61832 176936 61860
rect 151780 61820 151786 61832
rect 176930 61820 176936 61832
rect 176988 61820 176994 61872
rect 52362 61752 52368 61804
rect 52420 61792 52426 61804
rect 95786 61792 95792 61804
rect 52420 61764 95792 61792
rect 52420 61752 52426 61764
rect 95786 61752 95792 61764
rect 95844 61752 95850 61804
rect 97902 61752 97908 61804
rect 97960 61792 97966 61804
rect 133414 61792 133420 61804
rect 97960 61764 133420 61792
rect 97960 61752 97966 61764
rect 133414 61752 133420 61764
rect 133472 61752 133478 61804
rect 147582 61752 147588 61804
rect 147640 61792 147646 61804
rect 173986 61792 173992 61804
rect 147640 61764 173992 61792
rect 147640 61752 147646 61764
rect 173986 61752 173992 61764
rect 174044 61752 174050 61804
rect 18598 61684 18604 61736
rect 18656 61724 18662 61736
rect 54294 61724 54300 61736
rect 18656 61696 54300 61724
rect 18656 61684 18662 61696
rect 54294 61684 54300 61696
rect 54352 61684 54358 61736
rect 55122 61684 55128 61736
rect 55180 61724 55186 61736
rect 98546 61724 98552 61736
rect 55180 61696 98552 61724
rect 55180 61684 55186 61696
rect 98546 61684 98552 61696
rect 98604 61684 98610 61736
rect 140682 61684 140688 61736
rect 140740 61724 140746 61736
rect 168190 61724 168196 61736
rect 140740 61696 168196 61724
rect 140740 61684 140746 61696
rect 168190 61684 168196 61696
rect 168248 61684 168254 61736
rect 48222 61616 48228 61668
rect 48280 61656 48286 61668
rect 92842 61656 92848 61668
rect 48280 61628 92848 61656
rect 48280 61616 48286 61628
rect 92842 61616 92848 61628
rect 92900 61616 92906 61668
rect 95050 61616 95056 61668
rect 95108 61656 95114 61668
rect 130562 61656 130568 61668
rect 95108 61628 130568 61656
rect 95108 61616 95114 61628
rect 130562 61616 130568 61628
rect 130620 61616 130626 61668
rect 22002 61548 22008 61600
rect 22060 61588 22066 61600
rect 71590 61588 71596 61600
rect 22060 61560 71596 61588
rect 22060 61548 22066 61560
rect 71590 61548 71596 61560
rect 71648 61548 71654 61600
rect 77202 61548 77208 61600
rect 77260 61588 77266 61600
rect 116026 61588 116032 61600
rect 77260 61560 116032 61588
rect 77260 61548 77266 61560
rect 116026 61548 116032 61560
rect 116084 61548 116090 61600
rect 133230 61548 133236 61600
rect 133288 61588 133294 61600
rect 161474 61588 161480 61600
rect 133288 61560 161480 61588
rect 133288 61548 133294 61560
rect 161474 61548 161480 61560
rect 161532 61548 161538 61600
rect 17862 61480 17868 61532
rect 17920 61520 17926 61532
rect 67726 61520 67732 61532
rect 17920 61492 67732 61520
rect 17920 61480 17926 61492
rect 67726 61480 67732 61492
rect 67784 61480 67790 61532
rect 70302 61480 70308 61532
rect 70360 61520 70366 61532
rect 110230 61520 110236 61532
rect 70360 61492 110236 61520
rect 70360 61480 70366 61492
rect 110230 61480 110236 61492
rect 110288 61480 110294 61532
rect 131022 61480 131028 61532
rect 131080 61520 131086 61532
rect 160462 61520 160468 61532
rect 131080 61492 160468 61520
rect 131080 61480 131086 61492
rect 160462 61480 160468 61492
rect 160520 61480 160526 61532
rect 165522 61480 165528 61532
rect 165580 61520 165586 61532
rect 188522 61520 188528 61532
rect 165580 61492 188528 61520
rect 165580 61480 165586 61492
rect 188522 61480 188528 61492
rect 188580 61480 188586 61532
rect 517514 61480 517520 61532
rect 517572 61520 517578 61532
rect 564526 61520 564532 61532
rect 517572 61492 564532 61520
rect 517572 61480 517578 61492
rect 564526 61480 564532 61492
rect 564584 61480 564590 61532
rect 4890 61412 4896 61464
rect 4948 61452 4954 61464
rect 56134 61452 56140 61464
rect 4948 61424 56140 61452
rect 4948 61412 4954 61424
rect 56134 61412 56140 61424
rect 56192 61412 56198 61464
rect 73062 61412 73068 61464
rect 73120 61452 73126 61464
rect 113174 61452 113180 61464
rect 73120 61424 113180 61452
rect 73120 61412 73126 61424
rect 113174 61412 113180 61424
rect 113232 61412 113238 61464
rect 126882 61412 126888 61464
rect 126940 61452 126946 61464
rect 156506 61452 156512 61464
rect 126940 61424 156512 61452
rect 126940 61412 126946 61424
rect 156506 61412 156512 61424
rect 156564 61412 156570 61464
rect 162118 61412 162124 61464
rect 162176 61452 162182 61464
rect 185578 61452 185584 61464
rect 162176 61424 185584 61452
rect 162176 61412 162182 61424
rect 185578 61412 185584 61424
rect 185636 61412 185642 61464
rect 513098 61412 513104 61464
rect 513156 61452 513162 61464
rect 561674 61452 561680 61464
rect 513156 61424 561680 61452
rect 513156 61412 513162 61424
rect 561674 61412 561680 61424
rect 561732 61412 561738 61464
rect 8202 61344 8208 61396
rect 8260 61384 8266 61396
rect 59906 61384 59912 61396
rect 8260 61356 59912 61384
rect 8260 61344 8266 61356
rect 59906 61344 59912 61356
rect 59964 61344 59970 61396
rect 66162 61344 66168 61396
rect 66220 61384 66226 61396
rect 107378 61384 107384 61396
rect 66220 61356 107384 61384
rect 66220 61344 66226 61356
rect 107378 61344 107384 61356
rect 107436 61344 107442 61396
rect 111702 61344 111708 61396
rect 111760 61384 111766 61396
rect 144638 61384 144644 61396
rect 111760 61356 144644 61384
rect 111760 61344 111766 61356
rect 144638 61344 144644 61356
rect 144696 61344 144702 61396
rect 144730 61344 144736 61396
rect 144788 61384 144794 61396
rect 171134 61384 171140 61396
rect 144788 61356 171140 61384
rect 144788 61344 144794 61356
rect 171134 61344 171140 61356
rect 171192 61344 171198 61396
rect 173158 61344 173164 61396
rect 173216 61384 173222 61396
rect 194318 61384 194324 61396
rect 173216 61356 194324 61384
rect 173216 61344 173222 61356
rect 194318 61344 194324 61356
rect 194376 61344 194382 61396
rect 521746 61344 521752 61396
rect 521804 61384 521810 61396
rect 572806 61384 572812 61396
rect 521804 61356 572812 61384
rect 521804 61344 521810 61356
rect 572806 61344 572812 61356
rect 572864 61344 572870 61396
rect 130378 61276 130384 61328
rect 130436 61316 130442 61328
rect 157610 61316 157616 61328
rect 130436 61288 157616 61316
rect 130436 61276 130442 61288
rect 157610 61276 157616 61288
rect 157668 61276 157674 61328
rect 155218 61208 155224 61260
rect 155276 61248 155282 61260
rect 163406 61248 163412 61260
rect 155276 61220 163412 61248
rect 155276 61208 155282 61220
rect 163406 61208 163412 61220
rect 163464 61208 163470 61260
rect 533338 60664 533344 60716
rect 533396 60704 533402 60716
rect 580166 60704 580172 60716
rect 533396 60676 580172 60704
rect 533396 60664 533402 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2774 58896 2780 58948
rect 2832 58936 2838 58948
rect 4798 58936 4804 58948
rect 2832 58908 4804 58936
rect 2832 58896 2838 58908
rect 4798 58896 4804 58908
rect 4856 58896 4862 58948
rect 556798 46860 556804 46912
rect 556856 46900 556862 46912
rect 580166 46900 580172 46912
rect 556856 46872 580172 46900
rect 556856 46860 556862 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 33778 45540 33784 45552
rect 3568 45512 33784 45540
rect 3568 45500 3574 45512
rect 33778 45500 33784 45512
rect 33836 45500 33842 45552
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 29638 33096 29644 33108
rect 3568 33068 29644 33096
rect 3568 33056 3574 33068
rect 29638 33056 29644 33068
rect 29696 33056 29702 33108
rect 558178 33056 558184 33108
rect 558236 33096 558242 33108
rect 580166 33096 580172 33108
rect 558236 33068 580172 33096
rect 558236 33056 558242 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 511258 32376 511264 32428
rect 511316 32416 511322 32428
rect 557534 32416 557540 32428
rect 511316 32388 557540 32416
rect 511316 32376 511322 32388
rect 557534 32376 557540 32388
rect 557592 32376 557598 32428
rect 560938 20612 560944 20664
rect 560996 20652 561002 20664
rect 579982 20652 579988 20664
rect 560996 20624 579988 20652
rect 560996 20612 561002 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 292574 11704 292580 11756
rect 292632 11744 292638 11756
rect 293678 11744 293684 11756
rect 292632 11716 293684 11744
rect 292632 11704 292638 11716
rect 293678 11704 293684 11716
rect 293736 11704 293742 11756
rect 479518 8916 479524 8968
rect 479576 8956 479582 8968
rect 519538 8956 519544 8968
rect 479576 8928 519544 8956
rect 479576 8916 479582 8928
rect 519538 8916 519544 8928
rect 519596 8916 519602 8968
rect 520182 8916 520188 8968
rect 520240 8956 520246 8968
rect 569126 8956 569132 8968
rect 520240 8928 569132 8956
rect 520240 8916 520246 8928
rect 569126 8916 569132 8928
rect 569184 8916 569190 8968
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 35158 6848 35164 6860
rect 3476 6820 35164 6848
rect 3476 6808 3482 6820
rect 35158 6808 35164 6820
rect 35216 6808 35222 6860
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 86770 6196 86776 6248
rect 86828 6236 86834 6248
rect 124766 6236 124772 6248
rect 86828 6208 124772 6236
rect 86828 6196 86834 6208
rect 124766 6196 124772 6208
rect 124824 6196 124830 6248
rect 129366 6196 129372 6248
rect 129424 6236 129430 6248
rect 159542 6236 159548 6248
rect 129424 6208 159548 6236
rect 129424 6196 129430 6208
rect 159542 6196 159548 6208
rect 159600 6196 159606 6248
rect 58434 6128 58440 6180
rect 58492 6168 58498 6180
rect 101582 6168 101588 6180
rect 58492 6140 101588 6168
rect 58492 6128 58498 6140
rect 101582 6128 101588 6140
rect 101640 6128 101646 6180
rect 134610 6168 134616 6180
rect 103486 6140 134616 6168
rect 101030 6060 101036 6112
rect 101088 6100 101094 6112
rect 103486 6100 103514 6140
rect 134610 6128 134616 6140
rect 134668 6128 134674 6180
rect 169754 6128 169760 6180
rect 169812 6168 169818 6180
rect 191374 6168 191380 6180
rect 169812 6140 191380 6168
rect 169812 6128 169818 6140
rect 191374 6128 191380 6140
rect 191432 6128 191438 6180
rect 473262 6128 473268 6180
rect 473320 6168 473326 6180
rect 512454 6168 512460 6180
rect 473320 6140 512460 6168
rect 473320 6128 473326 6140
rect 512454 6128 512460 6140
rect 512512 6128 512518 6180
rect 101088 6072 103514 6100
rect 101088 6060 101094 6072
rect 472618 5448 472624 5500
rect 472676 5488 472682 5500
rect 508866 5488 508872 5500
rect 472676 5460 508872 5488
rect 472676 5448 472682 5460
rect 508866 5448 508872 5460
rect 508924 5448 508930 5500
rect 485130 5380 485136 5432
rect 485188 5420 485194 5432
rect 523034 5420 523040 5432
rect 485188 5392 523040 5420
rect 485188 5380 485194 5392
rect 523034 5380 523040 5392
rect 523092 5380 523098 5432
rect 410518 5312 410524 5364
rect 410576 5352 410582 5364
rect 434438 5352 434444 5364
rect 410576 5324 434444 5352
rect 410576 5312 410582 5324
rect 434438 5312 434444 5324
rect 434496 5312 434502 5364
rect 454678 5312 454684 5364
rect 454736 5352 454742 5364
rect 469858 5352 469864 5364
rect 454736 5324 469864 5352
rect 454736 5312 454742 5324
rect 469858 5312 469864 5324
rect 469916 5312 469922 5364
rect 476022 5312 476028 5364
rect 476080 5352 476086 5364
rect 515950 5352 515956 5364
rect 476080 5324 515956 5352
rect 476080 5312 476086 5324
rect 515950 5312 515956 5324
rect 516008 5312 516014 5364
rect 404170 5244 404176 5296
rect 404228 5284 404234 5296
rect 427262 5284 427268 5296
rect 404228 5256 427268 5284
rect 404228 5244 404234 5256
rect 427262 5244 427268 5256
rect 427320 5244 427326 5296
rect 433150 5244 433156 5296
rect 433208 5284 433214 5296
rect 462774 5284 462780 5296
rect 433208 5256 462780 5284
rect 433208 5244 433214 5256
rect 462774 5244 462780 5256
rect 462832 5244 462838 5296
rect 484302 5244 484308 5296
rect 484360 5284 484366 5296
rect 526622 5284 526628 5296
rect 484360 5256 526628 5284
rect 484360 5244 484366 5256
rect 526622 5244 526628 5256
rect 526680 5244 526686 5296
rect 383562 5176 383568 5228
rect 383620 5216 383626 5228
rect 402514 5216 402520 5228
rect 383620 5188 402520 5216
rect 383620 5176 383626 5188
rect 402514 5176 402520 5188
rect 402572 5176 402578 5228
rect 406930 5176 406936 5228
rect 406988 5216 406994 5228
rect 430850 5216 430856 5228
rect 406988 5188 430856 5216
rect 406988 5176 406994 5188
rect 430850 5176 430856 5188
rect 430908 5176 430914 5228
rect 447042 5176 447048 5228
rect 447100 5216 447106 5228
rect 480530 5216 480536 5228
rect 447100 5188 480536 5216
rect 447100 5176 447106 5188
rect 480530 5176 480536 5188
rect 480588 5176 480594 5228
rect 497550 5176 497556 5228
rect 497608 5216 497614 5228
rect 540790 5216 540796 5228
rect 497608 5188 540796 5216
rect 497608 5176 497614 5188
rect 540790 5176 540796 5188
rect 540848 5176 540854 5228
rect 386322 5108 386328 5160
rect 386380 5148 386386 5160
rect 406010 5148 406016 5160
rect 386380 5120 406016 5148
rect 386380 5108 386386 5120
rect 406010 5108 406016 5120
rect 406068 5108 406074 5160
rect 412542 5108 412548 5160
rect 412600 5148 412606 5160
rect 437934 5148 437940 5160
rect 412600 5120 437940 5148
rect 412600 5108 412606 5120
rect 437934 5108 437940 5120
rect 437992 5108 437998 5160
rect 453298 5108 453304 5160
rect 453356 5148 453362 5160
rect 487614 5148 487620 5160
rect 453356 5120 487620 5148
rect 453356 5108 453362 5120
rect 487614 5108 487620 5120
rect 487672 5108 487678 5160
rect 493962 5108 493968 5160
rect 494020 5148 494026 5160
rect 537202 5148 537208 5160
rect 494020 5120 537208 5148
rect 494020 5108 494026 5120
rect 537202 5108 537208 5120
rect 537260 5108 537266 5160
rect 389082 5040 389088 5092
rect 389140 5080 389146 5092
rect 409598 5080 409604 5092
rect 389140 5052 409604 5080
rect 389140 5040 389146 5052
rect 409598 5040 409604 5052
rect 409656 5040 409662 5092
rect 415302 5040 415308 5092
rect 415360 5080 415366 5092
rect 441430 5080 441436 5092
rect 415360 5052 441436 5080
rect 415360 5040 415366 5052
rect 441430 5040 441436 5052
rect 441488 5040 441494 5092
rect 449802 5040 449808 5092
rect 449860 5080 449866 5092
rect 484026 5080 484032 5092
rect 449860 5052 484032 5080
rect 449860 5040 449866 5052
rect 484026 5040 484032 5052
rect 484084 5040 484090 5092
rect 487062 5040 487068 5092
rect 487120 5080 487126 5092
rect 530118 5080 530124 5092
rect 487120 5052 530124 5080
rect 487120 5040 487126 5052
rect 530118 5040 530124 5052
rect 530176 5040 530182 5092
rect 392578 4972 392584 5024
rect 392636 5012 392642 5024
rect 413094 5012 413100 5024
rect 392636 4984 413100 5012
rect 392636 4972 392642 4984
rect 413094 4972 413100 4984
rect 413152 4972 413158 5024
rect 418062 4972 418068 5024
rect 418120 5012 418126 5024
rect 445018 5012 445024 5024
rect 418120 4984 445024 5012
rect 418120 4972 418126 4984
rect 445018 4972 445024 4984
rect 445076 4972 445082 5024
rect 455322 4972 455328 5024
rect 455380 5012 455386 5024
rect 491110 5012 491116 5024
rect 455380 4984 491116 5012
rect 455380 4972 455386 4984
rect 491110 4972 491116 4984
rect 491168 4972 491174 5024
rect 500218 4972 500224 5024
rect 500276 5012 500282 5024
rect 544286 5012 544292 5024
rect 500276 4984 544292 5012
rect 500276 4972 500282 4984
rect 544286 4972 544292 4984
rect 544344 4972 544350 5024
rect 394510 4904 394516 4956
rect 394568 4944 394574 4956
rect 416682 4944 416688 4956
rect 394568 4916 416688 4944
rect 394568 4904 394574 4916
rect 416682 4904 416688 4916
rect 416740 4904 416746 4956
rect 421558 4904 421564 4956
rect 421616 4944 421622 4956
rect 448606 4944 448612 4956
rect 421616 4916 448612 4944
rect 421616 4904 421622 4916
rect 448606 4904 448612 4916
rect 448664 4904 448670 4956
rect 458082 4904 458088 4956
rect 458140 4944 458146 4956
rect 494698 4944 494704 4956
rect 458140 4916 494704 4944
rect 458140 4904 458146 4916
rect 494698 4904 494704 4916
rect 494756 4904 494762 4956
rect 505002 4904 505008 4956
rect 505060 4944 505066 4956
rect 551462 4944 551468 4956
rect 505060 4916 551468 4944
rect 505060 4904 505066 4916
rect 551462 4904 551468 4916
rect 551520 4904 551526 4956
rect 62022 4836 62028 4888
rect 62080 4876 62086 4888
rect 104434 4876 104440 4888
rect 62080 4848 104440 4876
rect 62080 4836 62086 4848
rect 104434 4836 104440 4848
rect 104492 4836 104498 4888
rect 128354 4836 128360 4888
rect 128412 4876 128418 4888
rect 142154 4876 142160 4888
rect 128412 4848 142160 4876
rect 128412 4836 128418 4848
rect 142154 4836 142160 4848
rect 142212 4836 142218 4888
rect 397270 4836 397276 4888
rect 397328 4876 397334 4888
rect 420178 4876 420184 4888
rect 397328 4848 420184 4876
rect 397328 4836 397334 4848
rect 420178 4836 420184 4848
rect 420236 4836 420242 4888
rect 429010 4836 429016 4888
rect 429068 4876 429074 4888
rect 459186 4876 459192 4888
rect 429068 4848 459192 4876
rect 429068 4836 429074 4848
rect 459186 4836 459192 4848
rect 459244 4836 459250 4888
rect 462130 4836 462136 4888
rect 462188 4876 462194 4888
rect 498194 4876 498200 4888
rect 462188 4848 498200 4876
rect 462188 4836 462194 4848
rect 498194 4836 498200 4848
rect 498252 4836 498258 4888
rect 502242 4836 502248 4888
rect 502300 4876 502306 4888
rect 547874 4876 547880 4888
rect 502300 4848 547880 4876
rect 502300 4836 502306 4848
rect 547874 4836 547880 4848
rect 547932 4836 547938 4888
rect 30098 4768 30104 4820
rect 30156 4808 30162 4820
rect 72418 4808 72424 4820
rect 30156 4780 72424 4808
rect 30156 4768 30162 4780
rect 72418 4768 72424 4780
rect 72476 4768 72482 4820
rect 139394 4768 139400 4820
rect 139452 4808 139458 4820
rect 166258 4808 166264 4820
rect 139452 4780 166264 4808
rect 139452 4768 139458 4780
rect 166258 4768 166264 4780
rect 166316 4768 166322 4820
rect 381538 4768 381544 4820
rect 381596 4808 381602 4820
rect 398926 4808 398932 4820
rect 381596 4780 398932 4808
rect 381596 4768 381602 4780
rect 398926 4768 398932 4780
rect 398984 4768 398990 4820
rect 400030 4768 400036 4820
rect 400088 4808 400094 4820
rect 423766 4808 423772 4820
rect 400088 4780 423772 4808
rect 400088 4768 400094 4780
rect 423766 4768 423772 4780
rect 423824 4768 423830 4820
rect 426250 4768 426256 4820
rect 426308 4808 426314 4820
rect 455690 4808 455696 4820
rect 426308 4780 455696 4808
rect 426308 4768 426314 4780
rect 455690 4768 455696 4780
rect 455748 4768 455754 4820
rect 467742 4768 467748 4820
rect 467800 4808 467806 4820
rect 505370 4808 505376 4820
rect 467800 4780 505376 4808
rect 467800 4768 467806 4780
rect 505370 4768 505376 4780
rect 505428 4768 505434 4820
rect 507762 4768 507768 4820
rect 507820 4808 507826 4820
rect 554958 4808 554964 4820
rect 507820 4780 554964 4808
rect 507820 4768 507826 4780
rect 554958 4768 554964 4780
rect 555016 4768 555022 4820
rect 446398 4360 446404 4412
rect 446456 4400 446462 4412
rect 452102 4400 452108 4412
rect 446456 4372 452108 4400
rect 446456 4360 446462 4372
rect 452102 4360 452108 4372
rect 452160 4360 452166 4412
rect 442902 4156 442908 4208
rect 442960 4196 442966 4208
rect 442960 4168 446352 4196
rect 442960 4156 442966 4168
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 80698 4128 80704 4140
rect 45520 4100 80704 4128
rect 45520 4088 45526 4100
rect 80698 4088 80704 4100
rect 80756 4088 80762 4140
rect 108301 4131 108359 4137
rect 108301 4097 108313 4131
rect 108347 4128 108359 4131
rect 123386 4128 123392 4140
rect 108347 4100 123392 4128
rect 108347 4097 108359 4100
rect 108301 4091 108359 4097
rect 123386 4088 123392 4100
rect 123444 4088 123450 4140
rect 161290 4088 161296 4140
rect 161348 4128 161354 4140
rect 162118 4128 162124 4140
rect 161348 4100 162124 4128
rect 161348 4088 161354 4100
rect 162118 4088 162124 4100
rect 162176 4088 162182 4140
rect 322842 4088 322848 4140
rect 322900 4128 322906 4140
rect 327994 4128 328000 4140
rect 322900 4100 328000 4128
rect 322900 4088 322906 4100
rect 327994 4088 328000 4100
rect 328052 4088 328058 4140
rect 342162 4088 342168 4140
rect 342220 4128 342226 4140
rect 351638 4128 351644 4140
rect 342220 4100 351644 4128
rect 342220 4088 342226 4100
rect 351638 4088 351644 4100
rect 351696 4088 351702 4140
rect 355870 4088 355876 4140
rect 355928 4128 355934 4140
rect 368198 4128 368204 4140
rect 355928 4100 368204 4128
rect 355928 4088 355934 4100
rect 368198 4088 368204 4100
rect 368256 4088 368262 4140
rect 373902 4088 373908 4140
rect 373960 4128 373966 4140
rect 390646 4128 390652 4140
rect 373960 4100 390652 4128
rect 373960 4088 373966 4100
rect 390646 4088 390652 4100
rect 390704 4088 390710 4140
rect 397362 4088 397368 4140
rect 397420 4128 397426 4140
rect 418982 4128 418988 4140
rect 397420 4100 418988 4128
rect 397420 4088 397426 4100
rect 418982 4088 418988 4100
rect 419040 4088 419046 4140
rect 419442 4088 419448 4140
rect 419500 4128 419506 4140
rect 446214 4128 446220 4140
rect 419500 4100 446220 4128
rect 419500 4088 419506 4100
rect 446214 4088 446220 4100
rect 446272 4088 446278 4140
rect 446324 4128 446352 4168
rect 500310 4156 500316 4208
rect 500368 4196 500374 4208
rect 501782 4196 501788 4208
rect 500368 4168 501788 4196
rect 500368 4156 500374 4168
rect 501782 4156 501788 4168
rect 501840 4156 501846 4208
rect 529198 4156 529204 4208
rect 529256 4196 529262 4208
rect 533706 4196 533712 4208
rect 529256 4168 533712 4196
rect 529256 4156 529262 4168
rect 533706 4156 533712 4168
rect 533764 4156 533770 4208
rect 451093 4131 451151 4137
rect 451093 4128 451105 4131
rect 446324 4100 451105 4128
rect 451093 4097 451105 4100
rect 451139 4097 451151 4131
rect 451093 4091 451151 4097
rect 451182 4088 451188 4140
rect 451240 4128 451246 4140
rect 485222 4128 485228 4140
rect 451240 4100 485228 4128
rect 451240 4088 451246 4100
rect 485222 4088 485228 4100
rect 485280 4088 485286 4140
rect 487798 4088 487804 4140
rect 487856 4128 487862 4140
rect 507670 4128 507676 4140
rect 487856 4100 507676 4128
rect 487856 4088 487862 4100
rect 507670 4088 507676 4100
rect 507728 4088 507734 4140
rect 511902 4088 511908 4140
rect 511960 4128 511966 4140
rect 559742 4128 559748 4140
rect 511960 4100 559748 4128
rect 511960 4088 511966 4100
rect 559742 4088 559748 4100
rect 559800 4088 559806 4140
rect 31294 4020 31300 4072
rect 31352 4060 31358 4072
rect 43438 4060 43444 4072
rect 31352 4032 43444 4060
rect 31352 4020 31358 4032
rect 43438 4020 43444 4032
rect 43496 4020 43502 4072
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 90266 4060 90272 4072
rect 53800 4032 90272 4060
rect 53800 4020 53806 4032
rect 90266 4020 90272 4032
rect 90324 4020 90330 4072
rect 96246 4020 96252 4072
rect 96304 4060 96310 4072
rect 120718 4060 120724 4072
rect 96304 4032 120724 4060
rect 96304 4020 96310 4032
rect 120718 4020 120724 4032
rect 120776 4020 120782 4072
rect 344922 4020 344928 4072
rect 344980 4060 344986 4072
rect 355226 4060 355232 4072
rect 344980 4032 355232 4060
rect 344980 4020 344986 4032
rect 355226 4020 355232 4032
rect 355284 4020 355290 4072
rect 358722 4020 358728 4072
rect 358780 4060 358786 4072
rect 371694 4060 371700 4072
rect 358780 4032 371700 4060
rect 358780 4020 358786 4032
rect 371694 4020 371700 4032
rect 371752 4020 371758 4072
rect 375190 4020 375196 4072
rect 375248 4060 375254 4072
rect 393038 4060 393044 4072
rect 375248 4032 393044 4060
rect 375248 4020 375254 4032
rect 393038 4020 393044 4032
rect 393096 4020 393102 4072
rect 394602 4020 394608 4072
rect 394660 4060 394666 4072
rect 415486 4060 415492 4072
rect 394660 4032 415492 4060
rect 394660 4020 394666 4032
rect 415486 4020 415492 4032
rect 415544 4020 415550 4072
rect 422202 4020 422208 4072
rect 422260 4060 422266 4072
rect 449802 4060 449808 4072
rect 422260 4032 449808 4060
rect 422260 4020 422266 4032
rect 449802 4020 449808 4032
rect 449860 4020 449866 4072
rect 452473 4063 452531 4069
rect 452473 4029 452485 4063
rect 452519 4060 452531 4063
rect 456613 4063 456671 4069
rect 456613 4060 456625 4063
rect 452519 4032 456625 4060
rect 452519 4029 452531 4032
rect 452473 4023 452531 4029
rect 456613 4029 456625 4032
rect 456659 4029 456671 4063
rect 456613 4023 456671 4029
rect 456702 4020 456708 4072
rect 456760 4060 456766 4072
rect 492306 4060 492312 4072
rect 456760 4032 492312 4060
rect 456760 4020 456766 4032
rect 492306 4020 492312 4032
rect 492364 4020 492370 4072
rect 509142 4020 509148 4072
rect 509200 4060 509206 4072
rect 556154 4060 556160 4072
rect 509200 4032 556160 4060
rect 509200 4020 509206 4032
rect 556154 4020 556160 4032
rect 556212 4020 556218 4072
rect 41874 3952 41880 4004
rect 41932 3992 41938 4004
rect 79318 3992 79324 4004
rect 41932 3964 79324 3992
rect 41932 3952 41938 3964
rect 79318 3952 79324 3964
rect 79376 3952 79382 4004
rect 89162 3952 89168 4004
rect 89220 3992 89226 4004
rect 113818 3992 113824 4004
rect 89220 3964 113824 3992
rect 89220 3952 89226 3964
rect 113818 3952 113824 3964
rect 113876 3952 113882 4004
rect 128170 3952 128176 4004
rect 128228 3992 128234 4004
rect 146938 3992 146944 4004
rect 128228 3964 146944 3992
rect 128228 3952 128234 3964
rect 146938 3952 146944 3964
rect 146996 3952 147002 4004
rect 334618 3952 334624 4004
rect 334676 3992 334682 4004
rect 342162 3992 342168 4004
rect 334676 3964 342168 3992
rect 334676 3952 334682 3964
rect 342162 3952 342168 3964
rect 342220 3952 342226 4004
rect 343542 3952 343548 4004
rect 343600 3992 343606 4004
rect 354030 3992 354036 4004
rect 343600 3964 354036 3992
rect 343600 3952 343606 3964
rect 354030 3952 354036 3964
rect 354088 3952 354094 4004
rect 355962 3952 355968 4004
rect 356020 3992 356026 4004
rect 369394 3992 369400 4004
rect 356020 3964 369400 3992
rect 356020 3952 356026 3964
rect 369394 3952 369400 3964
rect 369452 3952 369458 4004
rect 372522 3952 372528 4004
rect 372580 3992 372586 4004
rect 389450 3992 389456 4004
rect 372580 3964 389456 3992
rect 372580 3952 372586 3964
rect 389450 3952 389456 3964
rect 389508 3952 389514 4004
rect 390278 3952 390284 4004
rect 390336 3992 390342 4004
rect 410794 3992 410800 4004
rect 390336 3964 410800 3992
rect 390336 3952 390342 3964
rect 410794 3952 410800 3964
rect 410852 3952 410858 4004
rect 413922 3952 413928 4004
rect 413980 3992 413986 4004
rect 439409 3995 439467 4001
rect 439409 3992 439421 3995
rect 413980 3964 439421 3992
rect 413980 3952 413986 3964
rect 439409 3961 439421 3964
rect 439455 3961 439467 3995
rect 439409 3955 439467 3961
rect 439498 3952 439504 4004
rect 439556 3992 439562 4004
rect 439556 3964 452700 3992
rect 439556 3952 439562 3964
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 69661 3927 69719 3933
rect 69661 3924 69673 3927
rect 38436 3896 69673 3924
rect 38436 3884 38442 3896
rect 69661 3893 69673 3896
rect 69707 3893 69719 3927
rect 69661 3887 69719 3893
rect 77386 3884 77392 3936
rect 77444 3924 77450 3936
rect 98641 3927 98699 3933
rect 98641 3924 98653 3927
rect 77444 3896 98653 3924
rect 77444 3884 77450 3896
rect 98641 3893 98653 3896
rect 98687 3893 98699 3927
rect 98641 3887 98699 3893
rect 99834 3884 99840 3936
rect 99892 3924 99898 3936
rect 108301 3927 108359 3933
rect 108301 3924 108313 3927
rect 99892 3896 108313 3924
rect 99892 3884 99898 3896
rect 108301 3893 108313 3896
rect 108347 3893 108359 3927
rect 128354 3924 128360 3936
rect 108301 3887 108359 3893
rect 108408 3896 128360 3924
rect 12250 3816 12256 3868
rect 12308 3856 12314 3868
rect 29730 3856 29736 3868
rect 12308 3828 29736 3856
rect 12308 3816 12314 3828
rect 29730 3816 29736 3828
rect 29788 3816 29794 3868
rect 34790 3816 34796 3868
rect 34848 3856 34854 3868
rect 75178 3856 75184 3868
rect 34848 3828 75184 3856
rect 34848 3816 34854 3828
rect 75178 3816 75184 3828
rect 75236 3816 75242 3868
rect 78582 3816 78588 3868
rect 78640 3856 78646 3868
rect 78640 3828 105952 3856
rect 78640 3816 78646 3828
rect 20530 3748 20536 3800
rect 20588 3788 20594 3800
rect 62758 3788 62764 3800
rect 20588 3760 62764 3788
rect 20588 3748 20594 3760
rect 62758 3748 62764 3760
rect 62816 3748 62822 3800
rect 65521 3791 65579 3797
rect 64846 3760 65472 3788
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 36538 3720 36544 3732
rect 1728 3692 36544 3720
rect 1728 3680 1734 3692
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 50982 3720 50988 3732
rect 50212 3692 50988 3720
rect 50212 3680 50218 3692
rect 50982 3680 50988 3692
rect 51040 3680 51046 3732
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 52362 3720 52368 3732
rect 51408 3692 52368 3720
rect 51408 3680 51414 3692
rect 52362 3680 52368 3692
rect 52420 3680 52426 3732
rect 52457 3723 52515 3729
rect 52457 3689 52469 3723
rect 52503 3720 52515 3723
rect 64846 3720 64874 3760
rect 52503 3692 64874 3720
rect 65444 3720 65472 3760
rect 65521 3757 65533 3791
rect 65567 3788 65579 3791
rect 69293 3791 69351 3797
rect 69293 3788 69305 3791
rect 65567 3760 69305 3788
rect 65567 3757 65579 3760
rect 65521 3751 65579 3757
rect 69293 3757 69305 3760
rect 69339 3757 69351 3791
rect 69293 3751 69351 3757
rect 69661 3791 69719 3797
rect 69661 3757 69673 3791
rect 69707 3788 69719 3791
rect 76558 3788 76564 3800
rect 69707 3760 76564 3788
rect 69707 3757 69719 3760
rect 69661 3751 69719 3757
rect 76558 3748 76564 3760
rect 76616 3748 76622 3800
rect 79321 3791 79379 3797
rect 79321 3757 79333 3791
rect 79367 3788 79379 3791
rect 98641 3791 98699 3797
rect 79367 3760 93854 3788
rect 79367 3757 79379 3760
rect 79321 3751 79379 3757
rect 88978 3720 88984 3732
rect 65444 3692 88984 3720
rect 52503 3689 52515 3692
rect 52457 3683 52515 3689
rect 88978 3680 88984 3692
rect 89036 3680 89042 3732
rect 93826 3720 93854 3760
rect 98641 3757 98653 3791
rect 98687 3788 98699 3791
rect 105538 3788 105544 3800
rect 98687 3760 105544 3788
rect 98687 3757 98699 3760
rect 98641 3751 98699 3757
rect 105538 3748 105544 3760
rect 105596 3748 105602 3800
rect 105924 3788 105952 3828
rect 108114 3816 108120 3868
rect 108172 3856 108178 3868
rect 108408 3856 108436 3896
rect 128354 3884 128360 3896
rect 128412 3884 128418 3936
rect 349062 3884 349068 3936
rect 349120 3924 349126 3936
rect 359918 3924 359924 3936
rect 349120 3896 359924 3924
rect 349120 3884 349126 3896
rect 359918 3884 359924 3896
rect 359976 3884 359982 3936
rect 362862 3884 362868 3936
rect 362920 3924 362926 3936
rect 377674 3924 377680 3936
rect 362920 3896 377680 3924
rect 362920 3884 362926 3896
rect 377674 3884 377680 3896
rect 377732 3884 377738 3936
rect 379422 3884 379428 3936
rect 379480 3924 379486 3936
rect 397730 3924 397736 3936
rect 379480 3896 397736 3924
rect 379480 3884 379486 3896
rect 397730 3884 397736 3896
rect 397788 3884 397794 3936
rect 398742 3884 398748 3936
rect 398800 3924 398806 3936
rect 421374 3924 421380 3936
rect 398800 3896 421380 3924
rect 398800 3884 398806 3896
rect 421374 3884 421380 3896
rect 421432 3884 421438 3936
rect 426342 3884 426348 3936
rect 426400 3924 426406 3936
rect 452565 3927 452623 3933
rect 452565 3924 452577 3927
rect 426400 3896 452577 3924
rect 426400 3884 426406 3896
rect 452565 3893 452577 3896
rect 452611 3893 452623 3927
rect 452672 3924 452700 3964
rect 453942 3952 453948 4004
rect 454000 3992 454006 4004
rect 488810 3992 488816 4004
rect 454000 3964 488816 3992
rect 454000 3952 454006 3964
rect 488810 3952 488816 3964
rect 488868 3952 488874 4004
rect 513190 3952 513196 4004
rect 513248 3992 513254 4004
rect 560846 3992 560852 4004
rect 513248 3964 560852 3992
rect 513248 3952 513254 3964
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 465166 3924 465172 3936
rect 452672 3896 465172 3924
rect 452565 3887 452623 3893
rect 465166 3884 465172 3896
rect 465224 3884 465230 3936
rect 497090 3924 497096 3936
rect 465736 3896 497096 3924
rect 108172 3828 108436 3856
rect 108172 3816 108178 3828
rect 109310 3816 109316 3868
rect 109368 3856 109374 3868
rect 116578 3856 116584 3868
rect 109368 3828 116584 3856
rect 109368 3816 109374 3828
rect 116578 3816 116584 3828
rect 116636 3816 116642 3868
rect 117590 3816 117596 3868
rect 117648 3856 117654 3868
rect 137278 3856 137284 3868
rect 117648 3828 137284 3856
rect 117648 3816 117654 3828
rect 137278 3816 137284 3828
rect 137336 3816 137342 3868
rect 314562 3816 314568 3868
rect 314620 3856 314626 3868
rect 318518 3856 318524 3868
rect 314620 3828 318524 3856
rect 314620 3816 314626 3828
rect 318518 3816 318524 3828
rect 318576 3816 318582 3868
rect 336550 3816 336556 3868
rect 336608 3856 336614 3868
rect 344649 3859 344707 3865
rect 344649 3856 344661 3859
rect 336608 3828 344661 3856
rect 336608 3816 336614 3828
rect 344649 3825 344661 3828
rect 344695 3825 344707 3859
rect 344649 3819 344707 3825
rect 346210 3816 346216 3868
rect 346268 3856 346274 3868
rect 356330 3856 356336 3868
rect 346268 3828 356336 3856
rect 346268 3816 346274 3828
rect 356330 3816 356336 3828
rect 356388 3816 356394 3868
rect 360102 3816 360108 3868
rect 360160 3856 360166 3868
rect 374086 3856 374092 3868
rect 360160 3828 374092 3856
rect 360160 3816 360166 3828
rect 374086 3816 374092 3828
rect 374144 3816 374150 3868
rect 380802 3816 380808 3868
rect 380860 3856 380866 3868
rect 400030 3856 400036 3868
rect 380860 3828 400036 3856
rect 380860 3816 380866 3828
rect 400030 3816 400036 3828
rect 400088 3816 400094 3868
rect 400122 3816 400128 3868
rect 400180 3856 400186 3868
rect 422570 3856 422576 3868
rect 400180 3828 422576 3856
rect 400180 3816 400186 3828
rect 422570 3816 422576 3828
rect 422628 3816 422634 3868
rect 424962 3816 424968 3868
rect 425020 3856 425026 3868
rect 453298 3856 453304 3868
rect 425020 3828 453304 3856
rect 425020 3816 425026 3828
rect 453298 3816 453304 3828
rect 453356 3816 453362 3868
rect 456613 3859 456671 3865
rect 456613 3825 456625 3859
rect 456659 3856 456671 3859
rect 460382 3856 460388 3868
rect 456659 3828 460388 3856
rect 456659 3825 456671 3828
rect 456613 3819 456671 3825
rect 460382 3816 460388 3828
rect 460440 3816 460446 3868
rect 460842 3816 460848 3868
rect 460900 3856 460906 3868
rect 465736 3856 465764 3896
rect 497090 3884 497096 3896
rect 497148 3884 497154 3936
rect 514662 3884 514668 3936
rect 514720 3924 514726 3936
rect 563238 3924 563244 3936
rect 514720 3896 563244 3924
rect 514720 3884 514726 3896
rect 563238 3884 563244 3896
rect 563296 3884 563302 3936
rect 495894 3856 495900 3868
rect 460900 3828 465764 3856
rect 465828 3828 495900 3856
rect 460900 3816 460906 3828
rect 108298 3788 108304 3800
rect 105924 3760 108304 3788
rect 108298 3748 108304 3760
rect 108356 3748 108362 3800
rect 114002 3748 114008 3800
rect 114060 3788 114066 3800
rect 135898 3788 135904 3800
rect 114060 3760 135904 3788
rect 114060 3748 114066 3760
rect 135898 3748 135904 3760
rect 135956 3748 135962 3800
rect 335262 3748 335268 3800
rect 335320 3788 335326 3800
rect 343358 3788 343364 3800
rect 335320 3760 343364 3788
rect 335320 3748 335326 3760
rect 343358 3748 343364 3760
rect 343416 3748 343422 3800
rect 350350 3748 350356 3800
rect 350408 3788 350414 3800
rect 362310 3788 362316 3800
rect 350408 3760 362316 3788
rect 350408 3748 350414 3760
rect 362310 3748 362316 3760
rect 362368 3748 362374 3800
rect 367002 3748 367008 3800
rect 367060 3788 367066 3800
rect 382366 3788 382372 3800
rect 367060 3760 382372 3788
rect 367060 3748 367066 3760
rect 382366 3748 382372 3760
rect 382424 3748 382430 3800
rect 384850 3748 384856 3800
rect 384908 3788 384914 3800
rect 403618 3788 403624 3800
rect 384908 3760 403624 3788
rect 384908 3748 384914 3760
rect 403618 3748 403624 3760
rect 403676 3748 403682 3800
rect 404262 3748 404268 3800
rect 404320 3788 404326 3800
rect 428458 3788 428464 3800
rect 404320 3760 428464 3788
rect 404320 3748 404326 3760
rect 428458 3748 428464 3760
rect 428516 3748 428522 3800
rect 430482 3748 430488 3800
rect 430540 3788 430546 3800
rect 452473 3791 452531 3797
rect 452473 3788 452485 3791
rect 430540 3760 452485 3788
rect 430540 3748 430546 3760
rect 452473 3757 452485 3760
rect 452519 3757 452531 3791
rect 452473 3751 452531 3757
rect 452565 3791 452623 3797
rect 452565 3757 452577 3791
rect 452611 3788 452623 3791
rect 454494 3788 454500 3800
rect 452611 3760 454500 3788
rect 452611 3757 452623 3760
rect 452565 3751 452623 3757
rect 454494 3748 454500 3760
rect 454552 3748 454558 3800
rect 465828 3788 465856 3828
rect 495894 3816 495900 3828
rect 495952 3816 495958 3868
rect 497458 3816 497464 3868
rect 497516 3856 497522 3868
rect 502886 3856 502892 3868
rect 497516 3828 502892 3856
rect 497516 3816 497522 3828
rect 502886 3816 502892 3828
rect 502944 3816 502950 3868
rect 516042 3816 516048 3868
rect 516100 3856 516106 3868
rect 564434 3856 564440 3868
rect 516100 3828 564440 3856
rect 516100 3816 516106 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 462240 3760 465856 3788
rect 465905 3791 465963 3797
rect 100110 3720 100116 3732
rect 93826 3692 100116 3720
rect 100110 3680 100116 3692
rect 100168 3680 100174 3732
rect 103330 3680 103336 3732
rect 103388 3720 103394 3732
rect 128998 3720 129004 3732
rect 103388 3692 129004 3720
rect 103388 3680 103394 3692
rect 128998 3680 129004 3692
rect 129056 3680 129062 3732
rect 132954 3680 132960 3732
rect 133012 3720 133018 3732
rect 151078 3720 151084 3732
rect 133012 3692 151084 3720
rect 133012 3680 133018 3692
rect 151078 3680 151084 3692
rect 151136 3680 151142 3732
rect 320910 3680 320916 3732
rect 320968 3720 320974 3732
rect 325510 3720 325516 3732
rect 320968 3692 325516 3720
rect 320968 3680 320974 3692
rect 325510 3680 325516 3692
rect 325568 3680 325574 3732
rect 325602 3680 325608 3732
rect 325660 3720 325666 3732
rect 331582 3720 331588 3732
rect 325660 3692 331588 3720
rect 325660 3680 325666 3692
rect 331582 3680 331588 3692
rect 331640 3680 331646 3732
rect 332318 3680 332324 3732
rect 332376 3720 332382 3732
rect 339862 3720 339868 3732
rect 332376 3692 339868 3720
rect 332376 3680 332382 3692
rect 339862 3680 339868 3692
rect 339920 3680 339926 3732
rect 340782 3680 340788 3732
rect 340840 3720 340846 3732
rect 350442 3720 350448 3732
rect 340840 3692 350448 3720
rect 340840 3680 340846 3692
rect 350442 3680 350448 3692
rect 350500 3680 350506 3732
rect 353202 3680 353208 3732
rect 353260 3720 353266 3732
rect 365806 3720 365812 3732
rect 353260 3692 365812 3720
rect 353260 3680 353266 3692
rect 365806 3680 365812 3692
rect 365864 3680 365870 3732
rect 368382 3680 368388 3732
rect 368440 3720 368446 3732
rect 384758 3720 384764 3732
rect 368440 3692 384764 3720
rect 368440 3680 368446 3692
rect 384758 3680 384764 3692
rect 384816 3680 384822 3732
rect 387610 3680 387616 3732
rect 387668 3720 387674 3732
rect 407206 3720 407212 3732
rect 387668 3692 407212 3720
rect 387668 3680 387674 3692
rect 407206 3680 407212 3692
rect 407264 3680 407270 3732
rect 413830 3680 413836 3732
rect 413888 3720 413894 3732
rect 439130 3720 439136 3732
rect 413888 3692 439136 3720
rect 413888 3680 413894 3692
rect 439130 3680 439136 3692
rect 439188 3680 439194 3732
rect 440142 3680 440148 3732
rect 440200 3720 440206 3732
rect 462041 3723 462099 3729
rect 462041 3720 462053 3723
rect 440200 3692 462053 3720
rect 440200 3680 440206 3692
rect 462041 3689 462053 3692
rect 462087 3689 462099 3723
rect 462041 3683 462099 3689
rect 18598 3652 18604 3664
rect 6886 3624 18604 3652
rect 566 3544 572 3596
rect 624 3584 630 3596
rect 6886 3584 6914 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 34609 3655 34667 3661
rect 18708 3624 34560 3652
rect 624 3556 6914 3584
rect 624 3544 630 3556
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 8812 3556 12480 3584
rect 8812 3544 8818 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4890 3516 4896 3528
rect 2924 3488 4896 3516
rect 2924 3476 2930 3488
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12452 3516 12480 3556
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 16482 3584 16488 3596
rect 15988 3556 16488 3584
rect 15988 3544 15994 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17862 3584 17868 3596
rect 17092 3556 17868 3584
rect 17092 3544 17098 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18708 3584 18736 3624
rect 18288 3556 18736 3584
rect 18288 3544 18294 3556
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 20622 3584 20628 3596
rect 19484 3556 20628 3584
rect 19484 3544 19490 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 24762 3584 24768 3596
rect 24268 3556 24768 3584
rect 24268 3544 24274 3556
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34532 3584 34560 3624
rect 34609 3621 34621 3655
rect 34655 3652 34667 3655
rect 65337 3655 65395 3661
rect 65337 3652 65349 3655
rect 34655 3624 65349 3652
rect 34655 3621 34667 3624
rect 34609 3615 34667 3621
rect 65337 3621 65349 3624
rect 65383 3621 65395 3655
rect 68738 3652 68744 3664
rect 65337 3615 65395 3621
rect 65444 3624 68744 3652
rect 65444 3584 65472 3624
rect 68738 3612 68744 3624
rect 68796 3612 68802 3664
rect 69293 3655 69351 3661
rect 69293 3621 69305 3655
rect 69339 3652 69351 3655
rect 73798 3652 73804 3664
rect 69339 3624 73804 3652
rect 69339 3621 69351 3624
rect 69293 3615 69351 3621
rect 73798 3612 73804 3624
rect 73856 3612 73862 3664
rect 74994 3612 75000 3664
rect 75052 3652 75058 3664
rect 106918 3652 106924 3664
rect 75052 3624 106924 3652
rect 75052 3612 75058 3624
rect 106918 3612 106924 3624
rect 106976 3612 106982 3664
rect 110506 3612 110512 3664
rect 110564 3652 110570 3664
rect 134518 3652 134524 3664
rect 110564 3624 134524 3652
rect 110564 3612 110570 3624
rect 134518 3612 134524 3624
rect 134576 3612 134582 3664
rect 156598 3652 156604 3664
rect 155328 3624 156604 3652
rect 34532 3556 65472 3584
rect 65518 3544 65524 3596
rect 65576 3584 65582 3596
rect 66162 3584 66168 3596
rect 65576 3556 66168 3584
rect 65576 3544 65582 3556
rect 66162 3544 66168 3556
rect 66220 3544 66226 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70302 3584 70308 3596
rect 69164 3556 70308 3584
rect 69164 3544 69170 3556
rect 70302 3544 70308 3556
rect 70360 3544 70366 3596
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 73062 3584 73068 3596
rect 72660 3556 73068 3584
rect 72660 3544 72666 3556
rect 73062 3544 73068 3556
rect 73120 3544 73126 3596
rect 76190 3544 76196 3596
rect 76248 3584 76254 3596
rect 77202 3584 77208 3596
rect 76248 3556 77208 3584
rect 76248 3544 76254 3556
rect 77202 3544 77208 3556
rect 77260 3544 77266 3596
rect 80882 3544 80888 3596
rect 80940 3584 80946 3596
rect 81342 3584 81348 3596
rect 80940 3556 81348 3584
rect 80940 3544 80946 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 82078 3544 82084 3596
rect 82136 3584 82142 3596
rect 113910 3584 113916 3596
rect 82136 3556 113916 3584
rect 82136 3544 82142 3556
rect 113910 3544 113916 3556
rect 113968 3544 113974 3596
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 115842 3584 115848 3596
rect 115256 3556 115848 3584
rect 115256 3544 115262 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 117222 3584 117228 3596
rect 116452 3556 117228 3584
rect 116452 3544 116458 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 118786 3544 118792 3596
rect 118844 3584 118850 3596
rect 119798 3584 119804 3596
rect 118844 3556 119804 3584
rect 118844 3544 118850 3556
rect 119798 3544 119804 3556
rect 119856 3544 119862 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 122742 3584 122748 3596
rect 122340 3556 122748 3584
rect 122340 3544 122346 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 124674 3544 124680 3596
rect 124732 3584 124738 3596
rect 125502 3584 125508 3596
rect 124732 3556 125508 3584
rect 124732 3544 124738 3556
rect 125502 3544 125508 3556
rect 125560 3544 125566 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 126882 3584 126888 3596
rect 125928 3556 126888 3584
rect 125928 3544 125934 3556
rect 126882 3544 126888 3556
rect 126940 3544 126946 3596
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 130378 3584 130384 3596
rect 127032 3556 130384 3584
rect 127032 3544 127038 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 130562 3544 130568 3596
rect 130620 3584 130626 3596
rect 131022 3584 131028 3596
rect 130620 3556 131028 3584
rect 130620 3544 130626 3556
rect 131022 3544 131028 3556
rect 131080 3544 131086 3596
rect 134150 3544 134156 3596
rect 134208 3584 134214 3596
rect 155218 3584 155224 3596
rect 134208 3556 155224 3584
rect 134208 3544 134214 3556
rect 155218 3544 155224 3556
rect 155276 3544 155282 3596
rect 57149 3519 57207 3525
rect 57149 3516 57161 3519
rect 12452 3488 57161 3516
rect 57149 3485 57161 3488
rect 57195 3485 57207 3519
rect 57149 3479 57207 3485
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64380 3488 93992 3516
rect 64380 3476 64386 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 58066 3448 58072 3460
rect 5316 3420 58072 3448
rect 5316 3408 5322 3420
rect 58066 3408 58072 3420
rect 58124 3408 58130 3460
rect 60826 3408 60832 3460
rect 60884 3448 60890 3460
rect 93857 3451 93915 3457
rect 93857 3448 93869 3451
rect 60884 3420 93869 3448
rect 60884 3408 60890 3420
rect 93857 3417 93869 3420
rect 93903 3417 93915 3451
rect 93964 3448 93992 3488
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 103422 3516 103428 3528
rect 102284 3488 103428 3516
rect 102284 3476 102290 3488
rect 103422 3476 103428 3488
rect 103480 3476 103486 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 133138 3516 133144 3528
rect 106976 3488 133144 3516
rect 106976 3476 106982 3488
rect 133138 3476 133144 3488
rect 133196 3476 133202 3528
rect 137370 3516 137376 3528
rect 134904 3488 137376 3516
rect 97258 3448 97264 3460
rect 93964 3420 97264 3448
rect 93857 3411 93915 3417
rect 97258 3408 97264 3420
rect 97316 3408 97322 3460
rect 104526 3408 104532 3460
rect 104584 3448 104590 3460
rect 134904 3448 134932 3488
rect 137370 3476 137376 3488
rect 137428 3476 137434 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 155328 3516 155356 3624
rect 156598 3612 156604 3624
rect 156656 3612 156662 3664
rect 171962 3612 171968 3664
rect 172020 3652 172026 3664
rect 173158 3652 173164 3664
rect 172020 3624 173164 3652
rect 172020 3612 172026 3624
rect 173158 3612 173164 3624
rect 173216 3612 173222 3664
rect 324222 3612 324228 3664
rect 324280 3652 324286 3664
rect 330386 3652 330392 3664
rect 324280 3624 330392 3652
rect 324280 3612 324286 3624
rect 330386 3612 330392 3624
rect 330444 3612 330450 3664
rect 331122 3612 331128 3664
rect 331180 3652 331186 3664
rect 338666 3652 338672 3664
rect 331180 3624 338672 3652
rect 331180 3612 331186 3624
rect 338666 3612 338672 3624
rect 338724 3612 338730 3664
rect 339402 3612 339408 3664
rect 339460 3652 339466 3664
rect 348050 3652 348056 3664
rect 339460 3624 348056 3652
rect 339460 3612 339466 3624
rect 348050 3612 348056 3624
rect 348108 3612 348114 3664
rect 348970 3612 348976 3664
rect 349028 3652 349034 3664
rect 361114 3652 361120 3664
rect 349028 3624 361120 3652
rect 349028 3612 349034 3624
rect 361114 3612 361120 3624
rect 361172 3612 361178 3664
rect 361390 3612 361396 3664
rect 361448 3652 361454 3664
rect 376478 3652 376484 3664
rect 361448 3624 376484 3652
rect 361448 3612 361454 3624
rect 376478 3612 376484 3624
rect 376536 3612 376542 3664
rect 382182 3612 382188 3664
rect 382240 3652 382246 3664
rect 401318 3652 401324 3664
rect 382240 3624 401324 3652
rect 382240 3612 382246 3624
rect 401318 3612 401324 3624
rect 401376 3612 401382 3664
rect 402882 3612 402888 3664
rect 402940 3652 402946 3664
rect 426158 3652 426164 3664
rect 402940 3624 426164 3652
rect 402940 3612 402946 3624
rect 426158 3612 426164 3624
rect 426216 3612 426222 3664
rect 427722 3612 427728 3664
rect 427780 3652 427786 3664
rect 456886 3652 456892 3664
rect 427780 3624 456892 3652
rect 427780 3612 427786 3624
rect 456886 3612 456892 3624
rect 456944 3612 456950 3664
rect 459462 3612 459468 3664
rect 459520 3652 459526 3664
rect 462240 3652 462268 3760
rect 465905 3757 465917 3791
rect 465951 3788 465963 3791
rect 499390 3788 499396 3800
rect 465951 3760 499396 3788
rect 465951 3757 465963 3760
rect 465905 3751 465963 3757
rect 499390 3748 499396 3760
rect 499448 3748 499454 3800
rect 518802 3748 518808 3800
rect 518860 3788 518866 3800
rect 568022 3788 568028 3800
rect 518860 3760 568028 3788
rect 518860 3748 518866 3760
rect 568022 3748 568028 3760
rect 568080 3748 568086 3800
rect 462317 3723 462375 3729
rect 462317 3689 462329 3723
rect 462363 3720 462375 3723
rect 462363 3692 464476 3720
rect 462363 3689 462375 3692
rect 462317 3683 462375 3689
rect 459520 3624 462268 3652
rect 459520 3612 459526 3624
rect 462406 3612 462412 3664
rect 462464 3652 462470 3664
rect 464448 3652 464476 3692
rect 466362 3680 466368 3732
rect 466420 3720 466426 3732
rect 466420 3692 472020 3720
rect 466420 3680 466426 3692
rect 471992 3652 472020 3692
rect 476758 3680 476764 3732
rect 476816 3720 476822 3732
rect 513558 3720 513564 3732
rect 476816 3692 513564 3720
rect 476816 3680 476822 3692
rect 513558 3680 513564 3692
rect 513616 3680 513622 3732
rect 517422 3680 517428 3732
rect 517480 3720 517486 3732
rect 566826 3720 566832 3732
rect 517480 3692 566832 3720
rect 517480 3680 517486 3692
rect 566826 3680 566832 3692
rect 566884 3680 566890 3732
rect 502889 3655 502947 3661
rect 502889 3652 502901 3655
rect 462464 3624 464108 3652
rect 464448 3624 470594 3652
rect 471992 3624 502901 3652
rect 462464 3612 462470 3624
rect 300762 3544 300768 3596
rect 300820 3584 300826 3596
rect 301958 3584 301964 3596
rect 300820 3556 301964 3584
rect 300820 3544 300826 3556
rect 301958 3544 301964 3556
rect 302016 3544 302022 3596
rect 303522 3544 303528 3596
rect 303580 3584 303586 3596
rect 305546 3584 305552 3596
rect 303580 3556 305552 3584
rect 303580 3544 303586 3556
rect 305546 3544 305552 3556
rect 305604 3544 305610 3596
rect 310422 3544 310428 3596
rect 310480 3584 310486 3596
rect 313826 3584 313832 3596
rect 310480 3556 313832 3584
rect 310480 3544 310486 3556
rect 313826 3544 313832 3556
rect 313884 3544 313890 3596
rect 317322 3544 317328 3596
rect 317380 3584 317386 3596
rect 320910 3584 320916 3596
rect 317380 3556 320916 3584
rect 317380 3544 317386 3556
rect 320910 3544 320916 3556
rect 320968 3544 320974 3596
rect 336642 3544 336648 3596
rect 336700 3584 336706 3596
rect 344554 3584 344560 3596
rect 336700 3556 344560 3584
rect 336700 3544 336706 3556
rect 344554 3544 344560 3556
rect 344612 3544 344618 3596
rect 344649 3587 344707 3593
rect 344649 3553 344661 3587
rect 344695 3584 344707 3587
rect 345750 3584 345756 3596
rect 344695 3556 345756 3584
rect 344695 3553 344707 3556
rect 344649 3547 344707 3553
rect 345750 3544 345756 3556
rect 345808 3544 345814 3596
rect 346302 3544 346308 3596
rect 346360 3584 346366 3596
rect 357526 3584 357532 3596
rect 346360 3556 357532 3584
rect 346360 3544 346366 3556
rect 357526 3544 357532 3556
rect 357584 3544 357590 3596
rect 358630 3544 358636 3596
rect 358688 3584 358694 3596
rect 372890 3584 372896 3596
rect 358688 3556 372896 3584
rect 358688 3544 358694 3556
rect 372890 3544 372896 3556
rect 372948 3544 372954 3596
rect 377950 3544 377956 3596
rect 378008 3584 378014 3596
rect 396534 3584 396540 3596
rect 378008 3556 396540 3584
rect 378008 3544 378014 3556
rect 396534 3544 396540 3556
rect 396592 3544 396598 3596
rect 405642 3544 405648 3596
rect 405700 3584 405706 3596
rect 429654 3584 429660 3596
rect 405700 3556 429660 3584
rect 405700 3544 405706 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 433242 3544 433248 3596
rect 433300 3584 433306 3596
rect 463970 3584 463976 3596
rect 433300 3556 463976 3584
rect 433300 3544 433306 3556
rect 463970 3544 463976 3556
rect 464028 3544 464034 3596
rect 464080 3584 464108 3624
rect 465905 3587 465963 3593
rect 465905 3584 465917 3587
rect 464080 3556 465917 3584
rect 465905 3553 465917 3556
rect 465951 3553 465963 3587
rect 465905 3547 465963 3553
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 467558 3584 467564 3596
rect 467156 3556 467564 3584
rect 467156 3544 467162 3556
rect 467558 3544 467564 3556
rect 467616 3544 467622 3596
rect 470566 3584 470594 3624
rect 502889 3621 502901 3624
rect 502935 3621 502947 3655
rect 502889 3615 502947 3621
rect 502978 3612 502984 3664
rect 503036 3652 503042 3664
rect 506474 3652 506480 3664
rect 503036 3624 506480 3652
rect 503036 3612 503042 3624
rect 506474 3612 506480 3624
rect 506532 3612 506538 3664
rect 521562 3612 521568 3664
rect 521620 3652 521626 3664
rect 571518 3652 571524 3664
rect 521620 3624 571524 3652
rect 521620 3612 521626 3624
rect 571518 3612 571524 3624
rect 571576 3612 571582 3664
rect 472250 3584 472256 3596
rect 470566 3556 472256 3584
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 511258 3584 511264 3596
rect 472452 3556 511264 3584
rect 140792 3488 155356 3516
rect 104584 3420 134932 3448
rect 104584 3408 104590 3420
rect 135254 3408 135260 3460
rect 135312 3448 135318 3460
rect 140792 3448 140820 3488
rect 155402 3476 155408 3528
rect 155460 3516 155466 3528
rect 155862 3516 155868 3528
rect 155460 3488 155868 3516
rect 155460 3476 155466 3488
rect 155862 3476 155868 3488
rect 155920 3476 155926 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 157242 3516 157248 3528
rect 156656 3488 157248 3516
rect 156656 3476 156662 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 165522 3516 165528 3528
rect 164936 3488 165528 3516
rect 164936 3476 164942 3488
rect 165522 3476 165528 3488
rect 165580 3476 165586 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 167178 3476 167184 3528
rect 167236 3516 167242 3528
rect 168282 3516 168288 3528
rect 167236 3488 168288 3516
rect 167236 3476 167242 3488
rect 168282 3476 168288 3488
rect 168340 3476 168346 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 189718 3476 189724 3528
rect 189776 3516 189782 3528
rect 190362 3516 190368 3528
rect 189776 3488 190368 3516
rect 189776 3476 189782 3488
rect 190362 3476 190368 3488
rect 190420 3476 190426 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 197906 3476 197912 3528
rect 197964 3516 197970 3528
rect 198642 3516 198648 3528
rect 197964 3488 198648 3516
rect 197964 3476 197970 3488
rect 198642 3476 198648 3488
rect 198700 3476 198706 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 200298 3476 200304 3528
rect 200356 3516 200362 3528
rect 201402 3516 201408 3528
rect 200356 3488 201408 3516
rect 200356 3476 200362 3488
rect 201402 3476 201408 3488
rect 201460 3476 201466 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 207382 3476 207388 3528
rect 207440 3516 207446 3528
rect 208302 3516 208308 3528
rect 207440 3488 208308 3516
rect 207440 3476 207446 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 211062 3516 211068 3528
rect 209832 3488 211068 3516
rect 209832 3476 209838 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 218054 3476 218060 3528
rect 218112 3516 218118 3528
rect 219158 3516 219164 3528
rect 218112 3488 219164 3516
rect 218112 3476 218118 3488
rect 219158 3476 219164 3488
rect 219216 3476 219222 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 225138 3476 225144 3528
rect 225196 3516 225202 3528
rect 226242 3516 226248 3528
rect 225196 3488 226248 3516
rect 225196 3476 225202 3488
rect 226242 3476 226248 3488
rect 226300 3476 226306 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227438 3516 227444 3528
rect 226392 3488 227444 3516
rect 226392 3476 226398 3488
rect 227438 3476 227444 3488
rect 227496 3476 227502 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235718 3516 235724 3528
rect 234672 3488 235724 3516
rect 234672 3476 234678 3488
rect 235718 3476 235724 3488
rect 235776 3476 235782 3528
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240778 3516 240784 3528
rect 239364 3488 240784 3516
rect 239364 3476 239370 3488
rect 240778 3476 240784 3488
rect 240836 3476 240842 3528
rect 241698 3476 241704 3528
rect 241756 3516 241762 3528
rect 242802 3516 242808 3528
rect 241756 3488 242808 3516
rect 241756 3476 241762 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244182 3516 244188 3528
rect 242952 3488 244188 3516
rect 242952 3476 242958 3488
rect 244182 3476 244188 3488
rect 244240 3476 244246 3528
rect 246390 3476 246396 3528
rect 246448 3516 246454 3528
rect 246942 3516 246948 3528
rect 246448 3488 246948 3516
rect 246448 3476 246454 3488
rect 246942 3476 246948 3488
rect 247000 3476 247006 3528
rect 247586 3476 247592 3528
rect 247644 3516 247650 3528
rect 248322 3516 248328 3528
rect 247644 3488 248328 3516
rect 247644 3476 247650 3488
rect 248322 3476 248328 3488
rect 248380 3476 248386 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252462 3516 252468 3528
rect 251232 3488 252468 3516
rect 251232 3476 251238 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 259454 3476 259460 3528
rect 259512 3516 259518 3528
rect 260558 3516 260564 3528
rect 259512 3488 260564 3516
rect 259512 3476 259518 3488
rect 260558 3476 260564 3488
rect 260616 3476 260622 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 265342 3476 265348 3528
rect 265400 3516 265406 3528
rect 266998 3516 267004 3528
rect 265400 3488 267004 3516
rect 265400 3476 265406 3488
rect 266998 3476 267004 3488
rect 267056 3476 267062 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 269758 3516 269764 3528
rect 267792 3488 269764 3516
rect 267792 3476 267798 3488
rect 269758 3476 269764 3488
rect 269816 3476 269822 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 274818 3476 274824 3528
rect 274876 3516 274882 3528
rect 275922 3516 275928 3528
rect 274876 3488 275928 3516
rect 274876 3476 274882 3488
rect 275922 3476 275928 3488
rect 275980 3476 275986 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 277302 3516 277308 3528
rect 276072 3488 277308 3516
rect 276072 3476 276078 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281902 3476 281908 3528
rect 281960 3516 281966 3528
rect 282822 3516 282828 3528
rect 281960 3488 282828 3516
rect 281960 3476 281966 3488
rect 282822 3476 282828 3488
rect 282880 3476 282886 3528
rect 283098 3476 283104 3528
rect 283156 3516 283162 3528
rect 285122 3516 285128 3528
rect 283156 3488 285128 3516
rect 283156 3476 283162 3488
rect 285122 3476 285128 3488
rect 285180 3476 285186 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 291838 3516 291844 3528
rect 291436 3488 291844 3516
rect 291436 3476 291442 3488
rect 291838 3476 291844 3488
rect 291896 3476 291902 3528
rect 303338 3476 303344 3528
rect 303396 3516 303402 3528
rect 304350 3516 304356 3528
rect 303396 3488 304356 3516
rect 303396 3476 303402 3488
rect 304350 3476 304356 3488
rect 304408 3476 304414 3528
rect 307662 3476 307668 3528
rect 307720 3516 307726 3528
rect 309042 3516 309048 3528
rect 307720 3488 309048 3516
rect 307720 3476 307726 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 311434 3516 311440 3528
rect 309836 3488 311440 3516
rect 309836 3476 309842 3488
rect 311434 3476 311440 3488
rect 311492 3476 311498 3528
rect 311802 3476 311808 3528
rect 311860 3516 311866 3528
rect 315022 3516 315028 3528
rect 311860 3488 315028 3516
rect 311860 3476 311866 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 318058 3476 318064 3528
rect 318116 3516 318122 3528
rect 319714 3516 319720 3528
rect 318116 3488 319720 3516
rect 318116 3476 318122 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 331858 3476 331864 3528
rect 331916 3516 331922 3528
rect 332686 3516 332692 3528
rect 331916 3488 332692 3516
rect 331916 3476 331922 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 339310 3476 339316 3528
rect 339368 3516 339374 3528
rect 349246 3516 349252 3528
rect 339368 3488 349252 3516
rect 339368 3476 339374 3488
rect 349246 3476 349252 3488
rect 349304 3476 349310 3528
rect 352558 3476 352564 3528
rect 352616 3516 352622 3528
rect 364610 3516 364616 3528
rect 352616 3488 364616 3516
rect 352616 3476 352622 3488
rect 364610 3476 364616 3488
rect 364668 3476 364674 3528
rect 365530 3476 365536 3528
rect 365588 3516 365594 3528
rect 381170 3516 381176 3528
rect 365588 3488 381176 3516
rect 365588 3476 365594 3488
rect 381170 3476 381176 3488
rect 381228 3476 381234 3528
rect 384942 3476 384948 3528
rect 385000 3516 385006 3528
rect 404814 3516 404820 3528
rect 385000 3488 404820 3516
rect 385000 3476 385006 3488
rect 404814 3476 404820 3488
rect 404872 3476 404878 3528
rect 407022 3476 407028 3528
rect 407080 3516 407086 3528
rect 432046 3516 432052 3528
rect 407080 3488 432052 3516
rect 407080 3476 407086 3488
rect 432046 3476 432052 3488
rect 432104 3476 432110 3528
rect 438762 3476 438768 3528
rect 438820 3516 438826 3528
rect 471054 3516 471060 3528
rect 438820 3488 471060 3516
rect 438820 3476 438826 3488
rect 471054 3476 471060 3488
rect 471112 3476 471118 3528
rect 471882 3476 471888 3528
rect 471940 3516 471946 3528
rect 472452 3516 472480 3556
rect 511258 3544 511264 3556
rect 511316 3544 511322 3596
rect 514018 3544 514024 3596
rect 514076 3584 514082 3596
rect 517146 3584 517152 3596
rect 514076 3556 517152 3584
rect 514076 3544 514082 3556
rect 517146 3544 517152 3556
rect 517204 3544 517210 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 529014 3584 529020 3596
rect 525116 3556 529020 3584
rect 525116 3544 525122 3556
rect 529014 3544 529020 3556
rect 529072 3544 529078 3596
rect 532050 3544 532056 3596
rect 532108 3584 532114 3596
rect 534902 3584 534908 3596
rect 532108 3556 534908 3584
rect 532108 3544 532114 3556
rect 534902 3544 534908 3556
rect 534960 3544 534966 3596
rect 534997 3587 535055 3593
rect 534997 3553 535009 3587
rect 535043 3584 535055 3587
rect 573910 3584 573916 3596
rect 535043 3556 573916 3584
rect 535043 3553 535055 3556
rect 534997 3547 535055 3553
rect 573910 3544 573916 3556
rect 573968 3544 573974 3596
rect 471940 3488 472480 3516
rect 471940 3476 471946 3488
rect 473998 3476 474004 3528
rect 474056 3516 474062 3528
rect 475746 3516 475752 3528
rect 474056 3488 475752 3516
rect 474056 3476 474062 3488
rect 475746 3476 475752 3488
rect 475804 3476 475810 3528
rect 480162 3476 480168 3528
rect 480220 3516 480226 3528
rect 520734 3516 520740 3528
rect 480220 3488 520740 3516
rect 480220 3476 480226 3488
rect 520734 3476 520740 3488
rect 520792 3476 520798 3528
rect 527082 3476 527088 3528
rect 527140 3516 527146 3528
rect 578602 3516 578608 3528
rect 527140 3488 578608 3516
rect 527140 3476 527146 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 135312 3420 140820 3448
rect 135312 3408 135318 3420
rect 141234 3408 141240 3460
rect 141292 3448 141298 3460
rect 142062 3448 142068 3460
rect 141292 3420 142068 3448
rect 141292 3408 141298 3420
rect 142062 3408 142068 3420
rect 142120 3408 142126 3460
rect 142430 3408 142436 3460
rect 142488 3448 142494 3460
rect 143442 3448 143448 3460
rect 142488 3420 143448 3448
rect 142488 3408 142494 3420
rect 143442 3408 143448 3420
rect 143500 3408 143506 3460
rect 143534 3408 143540 3460
rect 143592 3448 143598 3460
rect 144638 3448 144644 3460
rect 143592 3420 144644 3448
rect 143592 3408 143598 3420
rect 144638 3408 144644 3420
rect 144696 3408 144702 3460
rect 147122 3408 147128 3460
rect 147180 3448 147186 3460
rect 147582 3448 147588 3460
rect 147180 3420 147588 3448
rect 147180 3408 147186 3420
rect 147582 3408 147588 3420
rect 147640 3408 147646 3460
rect 148318 3408 148324 3460
rect 148376 3448 148382 3460
rect 148962 3448 148968 3460
rect 148376 3420 148968 3448
rect 148376 3408 148382 3420
rect 148962 3408 148968 3420
rect 149020 3408 149026 3460
rect 149514 3408 149520 3460
rect 149572 3448 149578 3460
rect 150342 3448 150348 3460
rect 149572 3420 150348 3448
rect 149572 3408 149578 3420
rect 150342 3408 150348 3420
rect 150400 3408 150406 3460
rect 150618 3408 150624 3460
rect 150676 3448 150682 3460
rect 151722 3448 151728 3460
rect 150676 3420 151728 3448
rect 150676 3408 150682 3420
rect 151722 3408 151728 3420
rect 151780 3408 151786 3460
rect 240502 3408 240508 3460
rect 240560 3448 240566 3460
rect 241422 3448 241428 3460
rect 240560 3420 241428 3448
rect 240560 3408 240566 3420
rect 241422 3408 241428 3420
rect 241480 3408 241486 3460
rect 248782 3408 248788 3460
rect 248840 3448 248846 3460
rect 249702 3448 249708 3460
rect 248840 3420 249708 3448
rect 248840 3408 248846 3420
rect 249702 3408 249708 3420
rect 249760 3408 249766 3460
rect 254670 3408 254676 3460
rect 254728 3448 254734 3460
rect 255958 3448 255964 3460
rect 254728 3420 255964 3448
rect 254728 3408 254734 3420
rect 255958 3408 255964 3420
rect 256016 3408 256022 3460
rect 266538 3408 266544 3460
rect 266596 3448 266602 3460
rect 267642 3448 267648 3460
rect 266596 3420 267648 3448
rect 266596 3408 266602 3420
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 286594 3408 286600 3460
rect 286652 3448 286658 3460
rect 287974 3448 287980 3460
rect 286652 3420 287980 3448
rect 286652 3408 286658 3420
rect 287974 3408 287980 3420
rect 288032 3408 288038 3460
rect 304902 3408 304908 3460
rect 304960 3448 304966 3460
rect 306742 3448 306748 3460
rect 304960 3420 306748 3448
rect 304960 3408 304966 3420
rect 306742 3408 306748 3420
rect 306800 3408 306806 3460
rect 307570 3408 307576 3460
rect 307628 3448 307634 3460
rect 310238 3448 310244 3460
rect 307628 3420 310244 3448
rect 307628 3408 307634 3420
rect 310238 3408 310244 3420
rect 310296 3408 310302 3460
rect 322750 3408 322756 3460
rect 322808 3448 322814 3460
rect 329190 3448 329196 3460
rect 322808 3420 329196 3448
rect 322808 3408 322814 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 332502 3408 332508 3460
rect 332560 3448 332566 3460
rect 340966 3448 340972 3460
rect 332560 3420 340972 3448
rect 332560 3408 332566 3420
rect 340966 3408 340972 3420
rect 341024 3408 341030 3460
rect 342070 3408 342076 3460
rect 342128 3448 342134 3460
rect 352834 3448 352840 3460
rect 342128 3420 352840 3448
rect 342128 3408 342134 3420
rect 352834 3408 352840 3420
rect 352892 3408 352898 3460
rect 357342 3408 357348 3460
rect 357400 3448 357406 3460
rect 370590 3448 370596 3460
rect 357400 3420 370596 3448
rect 357400 3408 357406 3420
rect 370590 3408 370596 3420
rect 370648 3408 370654 3460
rect 371050 3408 371056 3460
rect 371108 3448 371114 3460
rect 388254 3448 388260 3460
rect 371108 3420 388260 3448
rect 371108 3408 371114 3420
rect 388254 3408 388260 3420
rect 388312 3408 388318 3460
rect 390462 3408 390468 3460
rect 390520 3448 390526 3460
rect 411898 3448 411904 3460
rect 390520 3420 411904 3448
rect 390520 3408 390526 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 419350 3408 419356 3460
rect 419408 3448 419414 3460
rect 447410 3448 447416 3460
rect 419408 3420 447416 3448
rect 419408 3408 419414 3420
rect 447410 3408 447416 3420
rect 447468 3408 447474 3460
rect 448238 3408 448244 3460
rect 448296 3448 448302 3460
rect 481726 3448 481732 3460
rect 448296 3420 481732 3448
rect 448296 3408 448302 3420
rect 481726 3408 481732 3420
rect 481784 3408 481790 3460
rect 485682 3408 485688 3460
rect 485740 3448 485746 3460
rect 527818 3448 527824 3460
rect 485740 3420 527824 3448
rect 485740 3408 485746 3420
rect 527818 3408 527824 3420
rect 527876 3408 527882 3460
rect 528462 3408 528468 3460
rect 528520 3448 528526 3460
rect 580994 3448 581000 3460
rect 528520 3420 581000 3448
rect 528520 3408 528526 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26142 3380 26148 3392
rect 25372 3352 26148 3380
rect 25372 3340 25378 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 34609 3383 34667 3389
rect 34609 3380 34621 3383
rect 27764 3352 34621 3380
rect 27764 3340 27770 3352
rect 34609 3349 34621 3352
rect 34655 3349 34667 3383
rect 34609 3343 34667 3349
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 77938 3380 77944 3392
rect 43128 3352 77944 3380
rect 43128 3340 43134 3352
rect 77938 3340 77944 3352
rect 77996 3340 78002 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 84102 3380 84108 3392
rect 83332 3352 84108 3380
rect 83332 3340 83338 3352
rect 84102 3340 84108 3352
rect 84160 3340 84166 3392
rect 85666 3340 85672 3392
rect 85724 3380 85730 3392
rect 86862 3380 86868 3392
rect 85724 3352 86868 3380
rect 85724 3340 85730 3352
rect 86862 3340 86868 3352
rect 86920 3340 86926 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91097 3383 91155 3389
rect 91097 3349 91109 3383
rect 91143 3380 91155 3383
rect 107010 3380 107016 3392
rect 91143 3352 107016 3380
rect 91143 3349 91155 3352
rect 91097 3343 91155 3349
rect 107010 3340 107016 3352
rect 107068 3340 107074 3392
rect 121086 3340 121092 3392
rect 121144 3380 121150 3392
rect 138658 3380 138664 3392
rect 121144 3352 138664 3380
rect 121144 3340 121150 3352
rect 138658 3340 138664 3352
rect 138716 3340 138722 3392
rect 145926 3340 145932 3392
rect 145984 3380 145990 3392
rect 160738 3380 160744 3392
rect 145984 3352 160744 3380
rect 145984 3340 145990 3352
rect 160738 3340 160744 3352
rect 160796 3340 160802 3392
rect 313918 3340 313924 3392
rect 313976 3380 313982 3392
rect 317322 3380 317328 3392
rect 313976 3352 317328 3380
rect 313976 3340 313982 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 351822 3340 351828 3392
rect 351880 3380 351886 3392
rect 363506 3380 363512 3392
rect 351880 3352 363512 3380
rect 351880 3340 351886 3352
rect 363506 3340 363512 3352
rect 363564 3340 363570 3392
rect 369762 3340 369768 3392
rect 369820 3380 369826 3392
rect 385954 3380 385960 3392
rect 369820 3352 385960 3380
rect 369820 3340 369826 3352
rect 385954 3340 385960 3352
rect 386012 3340 386018 3392
rect 387702 3340 387708 3392
rect 387760 3380 387766 3392
rect 408402 3380 408408 3392
rect 387760 3352 408408 3380
rect 387760 3340 387766 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 409782 3340 409788 3392
rect 409840 3380 409846 3392
rect 435542 3380 435548 3392
rect 409840 3352 435548 3380
rect 409840 3340 409846 3352
rect 435542 3340 435548 3352
rect 435600 3340 435606 3392
rect 439409 3383 439467 3389
rect 439409 3349 439421 3383
rect 439455 3380 439467 3383
rect 440326 3380 440332 3392
rect 439455 3352 440332 3380
rect 439455 3349 439467 3352
rect 439409 3343 439467 3349
rect 440326 3340 440332 3352
rect 440384 3340 440390 3392
rect 441522 3340 441528 3392
rect 441580 3380 441586 3392
rect 473446 3380 473452 3392
rect 441580 3352 473452 3380
rect 441580 3340 441586 3352
rect 473446 3340 473452 3352
rect 473504 3340 473510 3392
rect 482830 3380 482836 3392
rect 480226 3352 482836 3380
rect 28902 3272 28908 3324
rect 28960 3312 28966 3324
rect 57149 3315 57207 3321
rect 28960 3284 57100 3312
rect 28960 3272 28966 3284
rect 35986 3204 35992 3256
rect 36044 3244 36050 3256
rect 57072 3244 57100 3284
rect 57149 3281 57161 3315
rect 57195 3312 57207 3315
rect 59998 3312 60004 3324
rect 57195 3284 60004 3312
rect 57195 3281 57207 3284
rect 57149 3275 57207 3281
rect 59998 3272 60004 3284
rect 60056 3272 60062 3324
rect 70302 3272 70308 3324
rect 70360 3312 70366 3324
rect 95878 3312 95884 3324
rect 70360 3284 89116 3312
rect 70360 3272 70366 3284
rect 61378 3244 61384 3256
rect 36044 3216 57008 3244
rect 57072 3216 61384 3244
rect 36044 3204 36050 3216
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 35250 3176 35256 3188
rect 26568 3148 35256 3176
rect 26568 3136 26574 3148
rect 35250 3136 35256 3148
rect 35308 3136 35314 3188
rect 37182 3136 37188 3188
rect 37240 3176 37246 3188
rect 37240 3148 45554 3176
rect 37240 3136 37246 3148
rect 45526 3108 45554 3148
rect 48958 3136 48964 3188
rect 49016 3176 49022 3188
rect 53098 3176 53104 3188
rect 49016 3148 53104 3176
rect 49016 3136 49022 3148
rect 53098 3136 53104 3148
rect 53156 3136 53162 3188
rect 55858 3108 55864 3120
rect 45526 3080 55864 3108
rect 55858 3068 55864 3080
rect 55916 3068 55922 3120
rect 56980 3108 57008 3216
rect 61378 3204 61384 3216
rect 61436 3204 61442 3256
rect 64138 3244 64144 3256
rect 61488 3216 64144 3244
rect 61488 3108 61516 3216
rect 64138 3204 64144 3216
rect 64196 3204 64202 3256
rect 66714 3204 66720 3256
rect 66772 3244 66778 3256
rect 84381 3247 84439 3253
rect 84381 3244 84393 3247
rect 66772 3216 84393 3244
rect 66772 3204 66778 3216
rect 84381 3213 84393 3216
rect 84427 3213 84439 3247
rect 89088 3244 89116 3284
rect 91204 3284 95884 3312
rect 91204 3244 91232 3284
rect 95878 3272 95884 3284
rect 95936 3272 95942 3324
rect 123478 3272 123484 3324
rect 123536 3312 123542 3324
rect 124122 3312 124128 3324
rect 123536 3284 124128 3312
rect 123536 3272 123542 3284
rect 124122 3272 124128 3284
rect 124180 3272 124186 3324
rect 131758 3272 131764 3324
rect 131816 3312 131822 3324
rect 133230 3312 133236 3324
rect 131816 3284 133236 3312
rect 131816 3272 131822 3284
rect 133230 3272 133236 3284
rect 133288 3272 133294 3324
rect 138842 3272 138848 3324
rect 138900 3312 138906 3324
rect 139302 3312 139308 3324
rect 138900 3284 139308 3312
rect 138900 3272 138906 3284
rect 139302 3272 139308 3284
rect 139360 3272 139366 3324
rect 163682 3272 163688 3324
rect 163740 3312 163746 3324
rect 164142 3312 164148 3324
rect 163740 3284 164148 3312
rect 163740 3272 163746 3284
rect 164142 3272 164148 3284
rect 164200 3272 164206 3324
rect 184934 3272 184940 3324
rect 184992 3312 184998 3324
rect 188338 3312 188344 3324
rect 184992 3284 188344 3312
rect 184992 3272 184998 3284
rect 188338 3272 188344 3284
rect 188396 3272 188402 3324
rect 229830 3272 229836 3324
rect 229888 3312 229894 3324
rect 230382 3312 230388 3324
rect 229888 3284 230388 3312
rect 229888 3272 229894 3284
rect 230382 3272 230388 3284
rect 230440 3272 230446 3324
rect 238110 3272 238116 3324
rect 238168 3312 238174 3324
rect 238662 3312 238668 3324
rect 238168 3284 238668 3312
rect 238168 3272 238174 3284
rect 238662 3272 238668 3284
rect 238720 3272 238726 3324
rect 257062 3272 257068 3324
rect 257120 3312 257126 3324
rect 257982 3312 257988 3324
rect 257120 3284 257988 3312
rect 257120 3272 257126 3284
rect 257982 3272 257988 3284
rect 258040 3272 258046 3324
rect 261754 3272 261760 3324
rect 261812 3312 261818 3324
rect 267090 3312 267096 3324
rect 261812 3284 267096 3312
rect 261812 3272 261818 3284
rect 267090 3272 267096 3284
rect 267148 3272 267154 3324
rect 272426 3272 272432 3324
rect 272484 3312 272490 3324
rect 276382 3312 276388 3324
rect 272484 3284 276388 3312
rect 272484 3272 272490 3284
rect 276382 3272 276388 3284
rect 276440 3272 276446 3324
rect 279510 3272 279516 3324
rect 279568 3312 279574 3324
rect 280798 3312 280804 3324
rect 279568 3284 280804 3312
rect 279568 3272 279574 3284
rect 280798 3272 280804 3284
rect 280856 3272 280862 3324
rect 306282 3272 306288 3324
rect 306340 3312 306346 3324
rect 307938 3312 307944 3324
rect 306340 3284 307944 3312
rect 306340 3272 306346 3284
rect 307938 3272 307944 3284
rect 307996 3272 308002 3324
rect 321002 3272 321008 3324
rect 321060 3312 321066 3324
rect 324406 3312 324412 3324
rect 321060 3284 324412 3312
rect 321060 3272 321066 3284
rect 324406 3272 324412 3284
rect 324464 3272 324470 3324
rect 328362 3272 328368 3324
rect 328420 3312 328426 3324
rect 335078 3312 335084 3324
rect 328420 3284 335084 3312
rect 328420 3272 328426 3284
rect 335078 3272 335084 3284
rect 335136 3272 335142 3324
rect 347682 3272 347688 3324
rect 347740 3312 347746 3324
rect 358722 3312 358728 3324
rect 347740 3284 358728 3312
rect 347740 3272 347746 3284
rect 358722 3272 358728 3284
rect 358780 3272 358786 3324
rect 361482 3272 361488 3324
rect 361540 3312 361546 3324
rect 375282 3312 375288 3324
rect 361540 3284 375288 3312
rect 361540 3272 361546 3284
rect 375282 3272 375288 3284
rect 375340 3272 375346 3324
rect 391842 3312 391848 3324
rect 375392 3284 391848 3312
rect 89088 3216 91232 3244
rect 84381 3207 84439 3213
rect 92750 3204 92756 3256
rect 92808 3244 92814 3256
rect 93762 3244 93768 3256
rect 92808 3216 93768 3244
rect 92808 3204 92814 3216
rect 93762 3204 93768 3216
rect 93820 3204 93826 3256
rect 93857 3247 93915 3253
rect 93857 3213 93869 3247
rect 93903 3244 93915 3247
rect 100018 3244 100024 3256
rect 93903 3216 100024 3244
rect 93903 3213 93915 3216
rect 93857 3207 93915 3213
rect 100018 3204 100024 3216
rect 100076 3204 100082 3256
rect 136450 3204 136456 3256
rect 136508 3244 136514 3256
rect 141418 3244 141424 3256
rect 136508 3216 141424 3244
rect 136508 3204 136514 3216
rect 141418 3204 141424 3216
rect 141476 3204 141482 3256
rect 318702 3204 318708 3256
rect 318760 3244 318766 3256
rect 323302 3244 323308 3256
rect 318760 3216 323308 3244
rect 318760 3204 318766 3216
rect 323302 3204 323308 3216
rect 323360 3204 323366 3256
rect 354582 3204 354588 3256
rect 354640 3244 354646 3256
rect 367002 3244 367008 3256
rect 354640 3216 367008 3244
rect 354640 3204 354646 3216
rect 367002 3204 367008 3216
rect 367060 3204 367066 3256
rect 375190 3204 375196 3256
rect 375248 3244 375254 3256
rect 375392 3244 375420 3284
rect 391842 3272 391848 3284
rect 391900 3272 391906 3324
rect 393222 3272 393228 3324
rect 393280 3312 393286 3324
rect 414290 3312 414296 3324
rect 393280 3284 414296 3312
rect 393280 3272 393286 3284
rect 414290 3272 414296 3284
rect 414348 3272 414354 3324
rect 416590 3272 416596 3324
rect 416648 3312 416654 3324
rect 442626 3312 442632 3324
rect 416648 3284 442632 3312
rect 416648 3272 416654 3284
rect 442626 3272 442632 3284
rect 442684 3272 442690 3324
rect 444282 3272 444288 3324
rect 444340 3312 444346 3324
rect 444340 3284 446536 3312
rect 444340 3272 444346 3284
rect 375248 3216 375420 3244
rect 375248 3204 375254 3216
rect 376662 3204 376668 3256
rect 376720 3244 376726 3256
rect 394234 3244 394240 3256
rect 376720 3216 394240 3244
rect 376720 3204 376726 3216
rect 394234 3204 394240 3216
rect 394292 3204 394298 3256
rect 411162 3204 411168 3256
rect 411220 3244 411226 3256
rect 436738 3244 436744 3256
rect 411220 3216 436744 3244
rect 411220 3204 411226 3216
rect 436738 3204 436744 3216
rect 436796 3204 436802 3256
rect 446508 3244 446536 3284
rect 448422 3272 448428 3324
rect 448480 3312 448486 3324
rect 480226 3312 480254 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 495342 3340 495348 3392
rect 495400 3380 495406 3392
rect 539594 3380 539600 3392
rect 495400 3352 539600 3380
rect 495400 3340 495406 3352
rect 539594 3340 539600 3352
rect 539652 3340 539658 3392
rect 541618 3340 541624 3392
rect 541676 3380 541682 3392
rect 543182 3380 543188 3392
rect 541676 3352 543188 3380
rect 541676 3340 541682 3352
rect 543182 3340 543188 3352
rect 543240 3340 543246 3392
rect 544378 3340 544384 3392
rect 544436 3380 544442 3392
rect 546865 3383 546923 3389
rect 544436 3352 546816 3380
rect 544436 3340 544442 3352
rect 448480 3284 480254 3312
rect 448480 3272 448486 3284
rect 482278 3272 482284 3324
rect 482336 3312 482342 3324
rect 500586 3312 500592 3324
rect 482336 3284 500592 3312
rect 482336 3272 482342 3284
rect 500586 3272 500592 3284
rect 500644 3272 500650 3324
rect 502889 3315 502947 3321
rect 502889 3281 502901 3315
rect 502935 3312 502947 3315
rect 504174 3312 504180 3324
rect 502935 3284 504180 3312
rect 502935 3281 502947 3284
rect 502889 3275 502947 3281
rect 504174 3272 504180 3284
rect 504232 3272 504238 3324
rect 508498 3272 508504 3324
rect 508556 3312 508562 3324
rect 510062 3312 510068 3324
rect 508556 3284 510068 3312
rect 508556 3272 508562 3284
rect 510062 3272 510068 3284
rect 510120 3272 510126 3324
rect 514021 3315 514079 3321
rect 514021 3281 514033 3315
rect 514067 3312 514079 3315
rect 542909 3315 542967 3321
rect 542909 3312 542921 3315
rect 514067 3284 542921 3312
rect 514067 3281 514079 3284
rect 514021 3275 514079 3281
rect 542909 3281 542921 3284
rect 542955 3281 542967 3315
rect 542909 3275 542967 3281
rect 542998 3272 543004 3324
rect 543056 3312 543062 3324
rect 546678 3312 546684 3324
rect 543056 3284 546684 3312
rect 543056 3272 543062 3284
rect 546678 3272 546684 3284
rect 546736 3272 546742 3324
rect 546788 3312 546816 3352
rect 546865 3349 546877 3383
rect 546911 3380 546923 3383
rect 577406 3380 577412 3392
rect 546911 3352 577412 3380
rect 546911 3349 546923 3352
rect 546865 3343 546923 3349
rect 577406 3340 577412 3352
rect 577464 3340 577470 3392
rect 550266 3312 550272 3324
rect 546788 3284 550272 3312
rect 550266 3272 550272 3284
rect 550324 3272 550330 3324
rect 551278 3272 551284 3324
rect 551336 3312 551342 3324
rect 575106 3312 575112 3324
rect 551336 3284 575112 3312
rect 551336 3272 551342 3284
rect 575106 3272 575112 3284
rect 575164 3272 575170 3324
rect 476942 3244 476948 3256
rect 441586 3216 446444 3244
rect 446508 3216 476948 3244
rect 61565 3179 61623 3185
rect 61565 3145 61577 3179
rect 61611 3176 61623 3179
rect 84838 3176 84844 3188
rect 61611 3148 84844 3176
rect 61611 3145 61623 3148
rect 61565 3139 61623 3145
rect 84838 3136 84844 3148
rect 84896 3136 84902 3188
rect 91554 3136 91560 3188
rect 91612 3176 91618 3188
rect 112438 3176 112444 3188
rect 91612 3148 112444 3176
rect 91612 3136 91618 3148
rect 112438 3136 112444 3148
rect 112496 3136 112502 3188
rect 193214 3136 193220 3188
rect 193272 3176 193278 3188
rect 194318 3176 194324 3188
rect 193272 3148 194324 3176
rect 193272 3136 193278 3148
rect 194318 3136 194324 3148
rect 194376 3136 194382 3188
rect 216858 3136 216864 3188
rect 216916 3176 216922 3188
rect 217962 3176 217968 3188
rect 216916 3148 217968 3176
rect 216916 3136 216922 3148
rect 217962 3136 217968 3148
rect 218020 3136 218026 3188
rect 310330 3136 310336 3188
rect 310388 3176 310394 3188
rect 312630 3176 312636 3188
rect 310388 3148 312636 3176
rect 310388 3136 310394 3148
rect 312630 3136 312636 3148
rect 312688 3136 312694 3188
rect 317230 3136 317236 3188
rect 317288 3176 317294 3188
rect 322106 3176 322112 3188
rect 317288 3148 322112 3176
rect 317288 3136 317294 3148
rect 322106 3136 322112 3148
rect 322164 3136 322170 3188
rect 329650 3136 329656 3188
rect 329708 3176 329714 3188
rect 336274 3176 336280 3188
rect 329708 3148 336280 3176
rect 329708 3136 329714 3148
rect 336274 3136 336280 3148
rect 336332 3136 336338 3188
rect 378042 3136 378048 3188
rect 378100 3176 378106 3188
rect 395338 3176 395344 3188
rect 378100 3148 395344 3176
rect 378100 3136 378106 3148
rect 395338 3136 395344 3148
rect 395396 3136 395402 3188
rect 408310 3136 408316 3188
rect 408368 3176 408374 3188
rect 433242 3176 433248 3188
rect 408368 3148 433248 3176
rect 408368 3136 408374 3148
rect 433242 3136 433248 3148
rect 433300 3136 433306 3188
rect 436002 3136 436008 3188
rect 436060 3176 436066 3188
rect 441586 3176 441614 3216
rect 436060 3148 441614 3176
rect 446416 3176 446444 3216
rect 476942 3204 476948 3216
rect 477000 3204 477006 3256
rect 489822 3204 489828 3256
rect 489880 3244 489886 3256
rect 532510 3244 532516 3256
rect 489880 3216 532516 3244
rect 489880 3204 489886 3216
rect 532510 3204 532516 3216
rect 532568 3204 532574 3256
rect 533430 3204 533436 3256
rect 533488 3244 533494 3256
rect 538398 3244 538404 3256
rect 533488 3216 538404 3244
rect 533488 3204 533494 3216
rect 538398 3204 538404 3216
rect 538456 3204 538462 3256
rect 576302 3244 576308 3256
rect 542372 3216 576308 3244
rect 467466 3176 467472 3188
rect 446416 3148 467472 3176
rect 436060 3136 436066 3148
rect 467466 3136 467472 3148
rect 467524 3136 467530 3188
rect 467558 3136 467564 3188
rect 467616 3176 467622 3188
rect 486418 3176 486424 3188
rect 467616 3148 486424 3176
rect 467616 3136 467622 3148
rect 486418 3136 486424 3148
rect 486476 3136 486482 3188
rect 503622 3136 503628 3188
rect 503680 3176 503686 3188
rect 514021 3179 514079 3185
rect 514021 3176 514033 3179
rect 503680 3148 514033 3176
rect 503680 3136 503686 3148
rect 514021 3145 514033 3148
rect 514067 3145 514079 3179
rect 514021 3139 514079 3145
rect 518360 3148 518894 3176
rect 56980 3080 61516 3108
rect 63218 3068 63224 3120
rect 63276 3108 63282 3120
rect 87598 3108 87604 3120
rect 63276 3080 87604 3108
rect 63276 3068 63282 3080
rect 87598 3068 87604 3080
rect 87656 3068 87662 3120
rect 168374 3068 168380 3120
rect 168432 3108 168438 3120
rect 169754 3108 169760 3120
rect 168432 3080 169760 3108
rect 168432 3068 168438 3080
rect 169754 3068 169760 3080
rect 169812 3068 169818 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 222102 3108 222108 3120
rect 221608 3080 222108 3108
rect 221608 3068 221614 3080
rect 222102 3068 222108 3080
rect 222160 3068 222166 3120
rect 313182 3068 313188 3120
rect 313240 3108 313246 3120
rect 316218 3108 316224 3120
rect 313240 3080 316224 3108
rect 313240 3068 313246 3080
rect 316218 3068 316224 3080
rect 316276 3068 316282 3120
rect 340230 3068 340236 3120
rect 340288 3108 340294 3120
rect 346946 3108 346952 3120
rect 340288 3080 346952 3108
rect 340288 3068 340294 3080
rect 346946 3068 346952 3080
rect 347004 3068 347010 3120
rect 371142 3068 371148 3120
rect 371200 3108 371206 3120
rect 387150 3108 387156 3120
rect 371200 3080 387156 3108
rect 371200 3068 371206 3080
rect 387150 3068 387156 3080
rect 387208 3068 387214 3120
rect 401502 3068 401508 3120
rect 401560 3108 401566 3120
rect 424962 3108 424968 3120
rect 401560 3080 424968 3108
rect 401560 3068 401566 3080
rect 424962 3068 424968 3080
rect 425020 3068 425026 3120
rect 437382 3068 437388 3120
rect 437440 3108 437446 3120
rect 468662 3108 468668 3120
rect 437440 3080 468668 3108
rect 437440 3068 437446 3080
rect 468662 3068 468668 3080
rect 468720 3068 468726 3120
rect 468757 3111 468815 3117
rect 468757 3077 468769 3111
rect 468803 3108 468815 3111
rect 478138 3108 478144 3120
rect 468803 3080 478144 3108
rect 468803 3077 468815 3080
rect 468757 3071 468815 3077
rect 478138 3068 478144 3080
rect 478196 3068 478202 3120
rect 483658 3068 483664 3120
rect 483716 3108 483722 3120
rect 518360 3108 518388 3148
rect 483716 3080 518388 3108
rect 518866 3108 518894 3148
rect 522850 3136 522856 3188
rect 522908 3176 522914 3188
rect 534997 3179 535055 3185
rect 534997 3176 535009 3179
rect 522908 3148 535009 3176
rect 522908 3136 522914 3148
rect 534997 3145 535009 3148
rect 535043 3145 535055 3179
rect 534997 3139 535055 3145
rect 540330 3136 540336 3188
rect 540388 3176 540394 3188
rect 542265 3179 542323 3185
rect 542265 3176 542277 3179
rect 540388 3148 542277 3176
rect 540388 3136 540394 3148
rect 542265 3145 542277 3148
rect 542311 3145 542323 3179
rect 542265 3139 542323 3145
rect 521838 3108 521844 3120
rect 518866 3080 521844 3108
rect 483716 3068 483722 3080
rect 521838 3068 521844 3080
rect 521896 3068 521902 3120
rect 526438 3068 526444 3120
rect 526496 3108 526502 3120
rect 531314 3108 531320 3120
rect 526496 3080 531320 3108
rect 526496 3068 526502 3080
rect 531314 3068 531320 3080
rect 531372 3068 531378 3120
rect 531958 3068 531964 3120
rect 532016 3108 532022 3120
rect 542372 3108 542400 3216
rect 576302 3204 576308 3216
rect 576360 3204 576366 3256
rect 570322 3176 570328 3188
rect 532016 3080 542400 3108
rect 542464 3148 570328 3176
rect 532016 3068 532022 3080
rect 44266 3000 44272 3052
rect 44324 3040 44330 3052
rect 65426 3040 65432 3052
rect 44324 3012 65432 3040
rect 44324 3000 44330 3012
rect 65426 3000 65432 3012
rect 65484 3000 65490 3052
rect 67910 3000 67916 3052
rect 67968 3040 67974 3052
rect 67968 3012 69796 3040
rect 67968 3000 67974 3012
rect 46658 2932 46664 2984
rect 46716 2972 46722 2984
rect 52457 2975 52515 2981
rect 52457 2972 52469 2975
rect 46716 2944 52469 2972
rect 46716 2932 46722 2944
rect 52457 2941 52469 2944
rect 52503 2941 52515 2975
rect 52457 2935 52515 2941
rect 56042 2932 56048 2984
rect 56100 2972 56106 2984
rect 69768 2972 69796 3012
rect 73798 3000 73804 3052
rect 73856 3040 73862 3052
rect 98546 3040 98552 3052
rect 73856 3012 98552 3040
rect 73856 3000 73862 3012
rect 98546 3000 98552 3012
rect 98604 3000 98610 3052
rect 151814 3000 151820 3052
rect 151872 3040 151878 3052
rect 152918 3040 152924 3052
rect 151872 3012 152924 3040
rect 151872 3000 151878 3012
rect 152918 3000 152924 3012
rect 152976 3000 152982 3052
rect 196802 3000 196808 3052
rect 196860 3040 196866 3052
rect 197262 3040 197268 3052
rect 196860 3012 197268 3040
rect 196860 3000 196866 3012
rect 197262 3000 197268 3012
rect 197320 3000 197326 3052
rect 321462 3000 321468 3052
rect 321520 3040 321526 3052
rect 326798 3040 326804 3052
rect 321520 3012 326804 3040
rect 321520 3000 321526 3012
rect 326798 3000 326804 3012
rect 326856 3000 326862 3052
rect 329742 3000 329748 3052
rect 329800 3040 329806 3052
rect 337470 3040 337476 3052
rect 329800 3012 337476 3040
rect 329800 3000 329806 3012
rect 337470 3000 337476 3012
rect 337528 3000 337534 3052
rect 368290 3000 368296 3052
rect 368348 3040 368354 3052
rect 383562 3040 383568 3052
rect 368348 3012 383568 3040
rect 368348 3000 368354 3012
rect 383562 3000 383568 3012
rect 383620 3000 383626 3052
rect 395982 3000 395988 3052
rect 396040 3040 396046 3052
rect 417878 3040 417884 3052
rect 396040 3012 417884 3040
rect 396040 3000 396046 3012
rect 417878 3000 417884 3012
rect 417936 3000 417942 3052
rect 431218 3000 431224 3052
rect 431276 3040 431282 3052
rect 443822 3040 443828 3052
rect 431276 3012 443828 3040
rect 431276 3000 431282 3012
rect 443822 3000 443828 3012
rect 443880 3000 443886 3052
rect 449158 3000 449164 3052
rect 449216 3040 449222 3052
rect 451093 3043 451151 3049
rect 449216 3012 451044 3040
rect 449216 3000 449222 3012
rect 79321 2975 79379 2981
rect 79321 2972 79333 2975
rect 56100 2944 69704 2972
rect 69768 2944 79333 2972
rect 56100 2932 56106 2944
rect 52546 2864 52552 2916
rect 52604 2904 52610 2916
rect 66898 2904 66904 2916
rect 52604 2876 66904 2904
rect 52604 2864 52610 2876
rect 66898 2864 66904 2876
rect 66956 2864 66962 2916
rect 69676 2904 69704 2944
rect 79321 2941 79333 2944
rect 79367 2941 79379 2975
rect 79321 2935 79379 2941
rect 84381 2975 84439 2981
rect 84381 2941 84393 2975
rect 84427 2972 84439 2975
rect 91738 2972 91744 2984
rect 84427 2944 91744 2972
rect 84427 2941 84439 2944
rect 84381 2935 84439 2941
rect 91738 2932 91744 2944
rect 91796 2932 91802 2984
rect 284294 2932 284300 2984
rect 284352 2972 284358 2984
rect 286042 2972 286048 2984
rect 284352 2944 286048 2972
rect 284352 2932 284358 2944
rect 286042 2932 286048 2944
rect 286100 2932 286106 2984
rect 326982 2932 326988 2984
rect 327040 2972 327046 2984
rect 333882 2972 333888 2984
rect 327040 2944 333888 2972
rect 327040 2932 327046 2944
rect 333882 2932 333888 2944
rect 333940 2932 333946 2984
rect 365622 2932 365628 2984
rect 365680 2972 365686 2984
rect 379974 2972 379980 2984
rect 365680 2944 379980 2972
rect 365680 2932 365686 2944
rect 379974 2932 379980 2944
rect 380032 2932 380038 2984
rect 436830 2932 436836 2984
rect 436888 2972 436894 2984
rect 450906 2972 450912 2984
rect 436888 2944 450912 2972
rect 436888 2932 436894 2944
rect 450906 2932 450912 2944
rect 450964 2932 450970 2984
rect 451016 2972 451044 3012
rect 451093 3009 451105 3043
rect 451139 3040 451151 3043
rect 474550 3040 474556 3052
rect 451139 3012 474556 3040
rect 451139 3009 451151 3012
rect 451093 3003 451151 3009
rect 474550 3000 474556 3012
rect 474608 3000 474614 3052
rect 490558 3000 490564 3052
rect 490616 3040 490622 3052
rect 514754 3040 514760 3052
rect 490616 3012 514760 3040
rect 490616 3000 490622 3012
rect 514754 3000 514760 3012
rect 514812 3000 514818 3052
rect 515490 3000 515496 3052
rect 515548 3040 515554 3052
rect 518342 3040 518348 3052
rect 515548 3012 518348 3040
rect 515548 3000 515554 3012
rect 518342 3000 518348 3012
rect 518400 3000 518406 3052
rect 518437 3043 518495 3049
rect 518437 3009 518449 3043
rect 518483 3040 518495 3043
rect 525426 3040 525432 3052
rect 518483 3012 525432 3040
rect 518483 3009 518495 3012
rect 518437 3003 518495 3009
rect 525426 3000 525432 3012
rect 525484 3000 525490 3052
rect 534718 3000 534724 3052
rect 534776 3040 534782 3052
rect 542464 3040 542492 3148
rect 570322 3136 570328 3148
rect 570380 3136 570386 3188
rect 545758 3068 545764 3120
rect 545816 3108 545822 3120
rect 582190 3108 582196 3120
rect 545816 3080 582196 3108
rect 545816 3068 545822 3080
rect 582190 3068 582196 3080
rect 582248 3068 582254 3120
rect 534776 3012 542492 3040
rect 542541 3043 542599 3049
rect 534776 3000 534782 3012
rect 542541 3009 542553 3043
rect 542587 3040 542599 3043
rect 552658 3040 552664 3052
rect 542587 3012 552664 3040
rect 542587 3009 542599 3012
rect 542541 3003 542599 3009
rect 552658 3000 552664 3012
rect 552716 3000 552722 3052
rect 582377 3043 582435 3049
rect 582377 3009 582389 3043
rect 582423 3040 582435 3043
rect 583386 3040 583392 3052
rect 582423 3012 583392 3040
rect 582423 3009 582435 3012
rect 582377 3003 582435 3009
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 479334 2972 479340 2984
rect 451016 2944 479340 2972
rect 479334 2932 479340 2944
rect 479392 2932 479398 2984
rect 482922 2932 482928 2984
rect 482980 2972 482986 2984
rect 524230 2972 524236 2984
rect 482980 2944 524236 2972
rect 482980 2932 482986 2944
rect 524230 2932 524236 2944
rect 524288 2932 524294 2984
rect 537478 2932 537484 2984
rect 537536 2972 537542 2984
rect 541986 2972 541992 2984
rect 537536 2944 541992 2972
rect 537536 2932 537542 2944
rect 541986 2932 541992 2944
rect 542044 2932 542050 2984
rect 546865 2975 546923 2981
rect 546865 2972 546877 2975
rect 542096 2944 546877 2972
rect 75270 2904 75276 2916
rect 69676 2876 75276 2904
rect 75270 2864 75276 2876
rect 75328 2864 75334 2916
rect 84470 2864 84476 2916
rect 84528 2904 84534 2916
rect 91097 2907 91155 2913
rect 91097 2904 91109 2907
rect 84528 2876 91109 2904
rect 84528 2864 84534 2876
rect 91097 2873 91109 2876
rect 91143 2873 91155 2907
rect 91097 2867 91155 2873
rect 93946 2864 93952 2916
rect 94004 2904 94010 2916
rect 95050 2904 95056 2916
rect 94004 2876 95056 2904
rect 94004 2864 94010 2876
rect 95050 2864 95056 2876
rect 95108 2864 95114 2916
rect 287790 2864 287796 2916
rect 287848 2904 287854 2916
rect 288342 2904 288348 2916
rect 287848 2876 288348 2904
rect 287848 2864 287854 2876
rect 288342 2864 288348 2876
rect 288400 2864 288406 2916
rect 364242 2864 364248 2916
rect 364300 2904 364306 2916
rect 378870 2904 378876 2916
rect 364300 2876 378876 2904
rect 364300 2864 364306 2876
rect 378870 2864 378876 2876
rect 378928 2864 378934 2916
rect 431862 2864 431868 2916
rect 431920 2904 431926 2916
rect 461578 2904 461584 2916
rect 431920 2876 461584 2904
rect 431920 2864 431926 2876
rect 461578 2864 461584 2876
rect 461636 2864 461642 2916
rect 464338 2864 464344 2916
rect 464396 2904 464402 2916
rect 468757 2907 468815 2913
rect 468757 2904 468769 2907
rect 464396 2876 468769 2904
rect 464396 2864 464402 2876
rect 468757 2873 468769 2876
rect 468803 2873 468815 2907
rect 468757 2867 468815 2873
rect 471238 2864 471244 2916
rect 471296 2904 471302 2916
rect 493502 2904 493508 2916
rect 471296 2876 493508 2904
rect 471296 2864 471302 2876
rect 493502 2864 493508 2876
rect 493560 2864 493566 2916
rect 515398 2864 515404 2916
rect 515456 2904 515462 2916
rect 518437 2907 518495 2913
rect 518437 2904 518449 2907
rect 515456 2876 518449 2904
rect 515456 2864 515462 2876
rect 518437 2873 518449 2876
rect 518483 2873 518495 2907
rect 518437 2867 518495 2873
rect 540238 2864 540244 2916
rect 540296 2904 540302 2916
rect 542096 2904 542124 2944
rect 546865 2941 546877 2944
rect 546911 2941 546923 2975
rect 546865 2935 546923 2941
rect 548518 2932 548524 2984
rect 548576 2972 548582 2984
rect 557350 2972 557356 2984
rect 548576 2944 557356 2972
rect 548576 2932 548582 2944
rect 557350 2932 557356 2944
rect 557408 2932 557414 2984
rect 540296 2876 542124 2904
rect 542909 2907 542967 2913
rect 540296 2864 540302 2876
rect 542909 2873 542921 2907
rect 542955 2904 542967 2907
rect 549070 2904 549076 2916
rect 542955 2876 549076 2904
rect 542955 2873 542967 2876
rect 542909 2867 542967 2873
rect 549070 2864 549076 2876
rect 549128 2864 549134 2916
rect 59630 2796 59636 2848
rect 59688 2836 59694 2848
rect 61565 2839 61623 2845
rect 61565 2836 61577 2839
rect 59688 2808 61577 2836
rect 59688 2796 59694 2808
rect 61565 2805 61577 2808
rect 61611 2805 61623 2839
rect 61565 2799 61623 2805
rect 137646 2796 137652 2848
rect 137704 2836 137710 2848
rect 139394 2836 139400 2848
rect 137704 2808 139400 2836
rect 137704 2796 137710 2808
rect 139394 2796 139400 2808
rect 139452 2796 139458 2848
rect 429102 2796 429108 2848
rect 429160 2836 429166 2848
rect 458082 2836 458088 2848
rect 429160 2808 458088 2836
rect 429160 2796 429166 2808
rect 458082 2796 458088 2808
rect 458140 2796 458146 2848
rect 468478 2796 468484 2848
rect 468536 2836 468542 2848
rect 489914 2836 489920 2848
rect 468536 2808 489920 2836
rect 468536 2796 468542 2808
rect 489914 2796 489920 2808
rect 489972 2796 489978 2848
rect 538858 2796 538864 2848
rect 538916 2836 538922 2848
rect 545482 2836 545488 2848
rect 538916 2808 545488 2836
rect 538916 2796 538922 2808
rect 545482 2796 545488 2808
rect 545540 2796 545546 2848
rect 547138 2796 547144 2848
rect 547196 2836 547202 2848
rect 553762 2836 553768 2848
rect 547196 2808 553768 2836
rect 547196 2796 547202 2808
rect 553762 2796 553768 2808
rect 553820 2796 553826 2848
<< via1 >>
rect 154120 700952 154172 701004
rect 327080 700952 327132 701004
rect 137836 700884 137888 700936
rect 322940 700884 322992 700936
rect 260748 700816 260800 700868
rect 462320 700816 462372 700868
rect 264888 700748 264940 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 339500 700680 339552 700732
rect 72976 700612 73028 700664
rect 335360 700612 335412 700664
rect 342904 700612 342956 700664
rect 364984 700612 365036 700664
rect 248328 700544 248380 700596
rect 527180 700544 527232 700596
rect 105452 700476 105504 700528
rect 166264 700476 166316 700528
rect 235172 700476 235224 700528
rect 242164 700476 242216 700528
rect 252468 700476 252520 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 343640 700408 343692 700460
rect 24308 700340 24360 700392
rect 351920 700340 351972 700392
rect 8116 700272 8168 700324
rect 347872 700272 347924 700324
rect 349804 700272 349856 700324
rect 429844 700272 429896 700324
rect 457444 700272 457496 700324
rect 494796 700272 494848 700324
rect 526444 700272 526496 700324
rect 559656 700272 559708 700324
rect 277308 700204 277360 700256
rect 413652 700204 413704 700256
rect 273168 700136 273220 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 310520 700068 310572 700120
rect 218980 700000 219032 700052
rect 314660 700000 314712 700052
rect 289728 699932 289780 699984
rect 348792 699932 348844 699984
rect 285588 699864 285640 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 298100 699796 298152 699848
rect 283840 699728 283892 699780
rect 302240 699728 302292 699780
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235908 696940 235960 696992
rect 580172 696940 580224 696992
rect 240048 683204 240100 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 356060 683136 356112 683188
rect 231768 670760 231820 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 364340 670692 364392 670744
rect 242164 668584 242216 668636
rect 306380 668584 306432 668636
rect 3424 656888 3476 656940
rect 360200 656888 360252 656940
rect 256332 643696 256384 643748
rect 457444 643696 457496 643748
rect 222936 643084 222988 643136
rect 580172 643084 580224 643136
rect 293960 642676 294012 642728
rect 299480 642676 299532 642728
rect 281356 642608 281408 642660
rect 342904 642608 342956 642660
rect 268844 642540 268896 642592
rect 349804 642540 349856 642592
rect 171048 642472 171100 642524
rect 318984 642472 319036 642524
rect 166264 642404 166316 642456
rect 331496 642404 331548 642456
rect 243820 642336 243872 642388
rect 526444 642336 526496 642388
rect 32404 641656 32456 641708
rect 486056 641656 486108 641708
rect 176936 641588 176988 641640
rect 369860 641588 369912 641640
rect 43536 641520 43588 641572
rect 390008 641520 390060 641572
rect 189448 641452 189500 641504
rect 536104 641452 536156 641504
rect 214564 641384 214616 641436
rect 569316 641384 569368 641436
rect 139400 641316 139452 641368
rect 189080 641316 189132 641368
rect 202052 641316 202104 641368
rect 558276 641316 558328 641368
rect 50436 641248 50488 641300
rect 423404 641248 423456 641300
rect 53196 641180 53248 641232
rect 435916 641180 435968 641232
rect 168564 641112 168616 641164
rect 551376 641112 551428 641164
rect 14464 641044 14516 641096
rect 402520 641044 402572 641096
rect 415860 641044 415912 641096
rect 477684 641044 477736 641096
rect 172796 640976 172848 641028
rect 562324 640976 562376 641028
rect 40684 640908 40736 640960
rect 440148 640908 440200 640960
rect 15844 640840 15896 640892
rect 415032 640840 415084 640892
rect 435364 640840 435416 640892
rect 527824 640840 527876 640892
rect 50344 640772 50396 640824
rect 452660 640772 452712 640824
rect 143540 640704 143592 640756
rect 547236 640704 547288 640756
rect 51724 640636 51776 640688
rect 461032 640636 461084 640688
rect 118516 640568 118568 640620
rect 543004 640568 543056 640620
rect 105912 640500 105964 640552
rect 531964 640500 532016 640552
rect 53104 640432 53156 640484
rect 490196 640432 490248 640484
rect 18604 640364 18656 640416
rect 465172 640364 465224 640416
rect 164424 640296 164476 640348
rect 175924 640296 175976 640348
rect 218704 640228 218756 640280
rect 538956 640228 539008 640280
rect 206192 640160 206244 640212
rect 537576 640160 537628 640212
rect 193680 640092 193732 640144
rect 536196 640092 536248 640144
rect 181168 640024 181220 640076
rect 533436 640024 533488 640076
rect 7656 639956 7708 640008
rect 369124 639956 369176 640008
rect 369860 639956 369912 640008
rect 580448 639956 580500 640008
rect 11796 639888 11848 639940
rect 381636 639888 381688 639940
rect 14556 639820 14608 639872
rect 394148 639820 394200 639872
rect 15936 639752 15988 639804
rect 406660 639752 406712 639804
rect 156052 639684 156104 639736
rect 548616 639684 548668 639736
rect 17316 639616 17368 639668
rect 419264 639616 419316 639668
rect 18696 639548 18748 639600
rect 431776 639548 431828 639600
rect 131028 639480 131080 639532
rect 544476 639480 544528 639532
rect 21456 639412 21508 639464
rect 444288 639412 444340 639464
rect 22744 639344 22796 639396
rect 456800 639344 456852 639396
rect 93400 639276 93452 639328
rect 530584 639276 530636 639328
rect 25504 639208 25556 639260
rect 469312 639208 469364 639260
rect 36544 639140 36596 639192
rect 481916 639140 481968 639192
rect 39304 639072 39356 639124
rect 494428 639072 494480 639124
rect 47584 639004 47636 639056
rect 506940 639004 506992 639056
rect 80888 638936 80940 638988
rect 540244 638936 540296 638988
rect 227076 638868 227128 638920
rect 530676 638868 530728 638920
rect 189080 638800 189132 638852
rect 580264 638800 580316 638852
rect 40868 638732 40920 638784
rect 377496 638732 377548 638784
rect 175924 638664 175976 638716
rect 580356 638664 580408 638716
rect 3516 638596 3568 638648
rect 415860 638596 415912 638648
rect 160560 638528 160612 638580
rect 537484 638528 537536 638580
rect 152280 638460 152332 638512
rect 532056 638460 532108 638512
rect 43444 638392 43496 638444
rect 448060 638392 448112 638444
rect 135260 638324 135312 638376
rect 538864 638324 538916 638376
rect 17224 638256 17276 638308
rect 427268 638256 427320 638308
rect 473360 638299 473412 638308
rect 473360 638265 473369 638299
rect 473369 638265 473403 638299
rect 473403 638265 473412 638299
rect 473360 638256 473412 638265
rect 502524 638299 502576 638308
rect 502524 638265 502533 638299
rect 502533 638265 502567 638299
rect 502567 638265 502576 638299
rect 502524 638256 502576 638265
rect 523316 638299 523368 638308
rect 523316 638265 523325 638299
rect 523325 638265 523359 638299
rect 523359 638265 523368 638299
rect 523316 638256 523368 638265
rect 148048 638188 148100 638240
rect 565084 638188 565136 638240
rect 126888 638120 126940 638172
rect 544384 638120 544436 638172
rect 114468 638052 114520 638104
rect 547144 638052 547196 638104
rect 102048 637984 102100 638036
rect 548524 637984 548576 638036
rect 97908 637959 97960 637968
rect 97908 637925 97917 637959
rect 97917 637925 97951 637959
rect 97951 637925 97960 637959
rect 97908 637916 97960 637925
rect 110328 637916 110380 637968
rect 122748 637916 122800 637968
rect 576124 637916 576176 637968
rect 89536 637848 89588 637900
rect 551284 637848 551336 637900
rect 574744 637780 574796 637832
rect 7564 637712 7616 637764
rect 573364 637644 573416 637696
rect 21364 637576 21416 637628
rect 35164 636828 35216 636880
rect 3332 632272 3384 632324
rect 7656 632272 7708 632324
rect 530676 632000 530728 632052
rect 579712 632000 579764 632052
rect 3608 619556 3660 619608
rect 40868 619556 40920 619608
rect 538956 618196 539008 618248
rect 579804 618196 579856 618248
rect 3056 607112 3108 607164
rect 32496 607112 32548 607164
rect 565176 591948 565228 592000
rect 580172 591948 580224 592000
rect 3332 580932 3384 580984
rect 11796 580932 11848 580984
rect 569316 578144 569368 578196
rect 580172 578144 580224 578196
rect 3332 567128 3384 567180
rect 43536 567128 43588 567180
rect 537576 564340 537628 564392
rect 580172 564340 580224 564392
rect 3332 554684 3384 554736
rect 33876 554684 33928 554736
rect 562416 538160 562468 538212
rect 580172 538160 580224 538212
rect 3332 528504 3384 528556
rect 14556 528504 14608 528556
rect 558276 525716 558328 525768
rect 580172 525716 580224 525768
rect 3148 516060 3200 516112
rect 14464 516060 14516 516112
rect 536196 511912 536248 511964
rect 580172 511912 580224 511964
rect 2964 502256 3016 502308
rect 35256 502256 35308 502308
rect 561128 485732 561180 485784
rect 580172 485732 580224 485784
rect 3240 476008 3292 476060
rect 15936 476008 15988 476060
rect 536104 471928 536156 471980
rect 580172 471928 580224 471980
rect 3056 463632 3108 463684
rect 15844 463632 15896 463684
rect 533436 458124 533488 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 40776 449828 40828 449880
rect 562324 431876 562376 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 17316 423580 17368 423632
rect 2964 411204 3016 411256
rect 17224 411204 17276 411256
rect 551376 405628 551428 405680
rect 580172 405628 580224 405680
rect 3332 398760 3384 398812
rect 50436 398760 50488 398812
rect 537484 379448 537536 379500
rect 580172 379448 580224 379500
rect 3332 372512 3384 372564
rect 18696 372512 18748 372564
rect 3332 358708 3384 358760
rect 40684 358708 40736 358760
rect 548616 353200 548668 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 53196 346332 53248 346384
rect 565084 325592 565136 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 21456 320084 21508 320136
rect 532056 313216 532108 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 50344 306280 50396 306332
rect 547236 299412 547288 299464
rect 579620 299412 579672 299464
rect 3332 293904 3384 293956
rect 43444 293904 43496 293956
rect 538864 273164 538916 273216
rect 579896 273164 579948 273216
rect 2964 267656 3016 267708
rect 22744 267656 22796 267708
rect 3148 255212 3200 255264
rect 18604 255212 18656 255264
rect 544476 245556 544528 245608
rect 580172 245556 580224 245608
rect 3240 241408 3292 241460
rect 51724 241408 51776 241460
rect 576124 233180 576176 233232
rect 579988 233180 580040 233232
rect 544384 219376 544436 219428
rect 580172 219376 580224 219428
rect 3332 215228 3384 215280
rect 25504 215228 25556 215280
rect 543004 206932 543056 206984
rect 579804 206932 579856 206984
rect 574744 193128 574796 193180
rect 580172 193128 580224 193180
rect 3516 188844 3568 188896
rect 7564 188844 7616 188896
rect 547144 179324 547196 179376
rect 580172 179324 580224 179376
rect 531964 166948 532016 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 36544 164160 36596 164212
rect 573364 153144 573416 153196
rect 580172 153144 580224 153196
rect 3516 150356 3568 150408
rect 53104 150356 53156 150408
rect 548524 139340 548576 139392
rect 580172 139340 580224 139392
rect 3516 137912 3568 137964
rect 32404 137912 32456 137964
rect 530584 126896 530636 126948
rect 580172 126896 580224 126948
rect 569224 113092 569276 113144
rect 579804 113092 579856 113144
rect 3148 111732 3200 111784
rect 39304 111732 39356 111784
rect 551284 100648 551336 100700
rect 580172 100648 580224 100700
rect 3516 97928 3568 97980
rect 21364 97928 21416 97980
rect 540244 86912 540296 86964
rect 580172 86912 580224 86964
rect 3516 85484 3568 85536
rect 11704 85484 11756 85536
rect 566464 73108 566516 73160
rect 580172 73108 580224 73160
rect 3516 71680 3568 71732
rect 47584 71680 47636 71732
rect 23388 63452 23440 63504
rect 72608 63452 72660 63504
rect 84844 63452 84896 63504
rect 102508 63452 102560 63504
rect 105544 63452 105596 63504
rect 117044 63452 117096 63504
rect 119804 63452 119856 63504
rect 150808 63452 150860 63504
rect 157248 63452 157300 63504
rect 181720 63452 181772 63504
rect 183468 63452 183520 63504
rect 202972 63452 203024 63504
rect 209688 63452 209740 63504
rect 224224 63452 224276 63504
rect 229008 63452 229060 63504
rect 240692 63452 240744 63504
rect 248328 63452 248380 63504
rect 256148 63452 256200 63504
rect 499580 63452 499632 63504
rect 538864 63452 538916 63504
rect 24768 63384 24820 63436
rect 73528 63384 73580 63436
rect 87604 63384 87656 63436
rect 105452 63384 105504 63436
rect 115848 63384 115900 63436
rect 147956 63384 148008 63436
rect 153016 63384 153068 63436
rect 177856 63384 177908 63436
rect 186228 63384 186280 63436
rect 205916 63384 205968 63436
rect 211068 63384 211120 63436
rect 225236 63384 225288 63436
rect 226248 63384 226300 63436
rect 237748 63384 237800 63436
rect 240784 63384 240836 63436
rect 249340 63384 249392 63436
rect 470600 63384 470652 63436
rect 508504 63384 508556 63436
rect 509240 63384 509292 63436
rect 548524 63384 548576 63436
rect 26148 63316 26200 63368
rect 74540 63316 74592 63368
rect 75276 63316 75328 63368
rect 99656 63316 99708 63368
rect 106188 63316 106240 63368
rect 140228 63316 140280 63368
rect 148968 63316 149020 63368
rect 175004 63316 175056 63368
rect 177948 63316 178000 63368
rect 198188 63316 198240 63368
rect 198648 63316 198700 63368
rect 215576 63316 215628 63368
rect 219256 63316 219308 63368
rect 231952 63316 232004 63368
rect 233148 63316 233200 63368
rect 243544 63316 243596 63368
rect 244188 63316 244240 63368
rect 252284 63316 252336 63368
rect 334348 63316 334400 63368
rect 335268 63316 335320 63368
rect 353668 63316 353720 63368
rect 354588 63316 354640 63368
rect 372988 63316 373040 63368
rect 373908 63316 373960 63368
rect 392308 63316 392360 63368
rect 393228 63316 393280 63368
rect 411628 63316 411680 63368
rect 412548 63316 412600 63368
rect 445484 63316 445536 63368
rect 449164 63316 449216 63368
rect 457076 63316 457128 63368
rect 471244 63316 471296 63368
rect 494704 63316 494756 63368
rect 495348 63316 495400 63368
rect 20628 63248 20680 63300
rect 69664 63248 69716 63300
rect 79416 63248 79468 63300
rect 88064 63248 88116 63300
rect 90364 63248 90416 63300
rect 97724 63248 97776 63300
rect 99288 63248 99340 63300
rect 134432 63248 134484 63300
rect 138664 63248 138716 63300
rect 152740 63248 152792 63300
rect 154488 63248 154540 63300
rect 179788 63248 179840 63300
rect 180708 63248 180760 63300
rect 201040 63248 201092 63300
rect 204168 63248 204220 63300
rect 220360 63248 220412 63300
rect 223488 63248 223540 63300
rect 235816 63248 235868 63300
rect 235908 63248 235960 63300
rect 246488 63248 246540 63300
rect 454132 63248 454184 63300
rect 468484 63248 468536 63300
rect 482192 63248 482244 63300
rect 482928 63248 482980 63300
rect 493784 63248 493836 63300
rect 533436 63316 533488 63368
rect 496636 63248 496688 63300
rect 537484 63248 537536 63300
rect 10968 63180 11020 63232
rect 61936 63180 61988 63232
rect 77392 63180 77444 63232
rect 77944 63180 77996 63232
rect 88984 63180 89036 63232
rect 93768 63180 93820 63232
rect 129556 63180 129608 63232
rect 134524 63180 134576 63232
rect 144092 63180 144144 63232
rect 144828 63180 144880 63232
rect 172060 63180 172112 63232
rect 175188 63180 175240 63232
rect 196256 63180 196308 63232
rect 197268 63180 197320 63232
rect 214564 63180 214616 63232
rect 215208 63180 215260 63232
rect 229100 63180 229152 63232
rect 231768 63180 231820 63232
rect 242624 63180 242676 63232
rect 246948 63180 247000 63232
rect 255136 63180 255188 63232
rect 439688 63180 439740 63232
rect 440148 63180 440200 63232
rect 462872 63180 462924 63232
rect 482284 63180 482336 63232
rect 489920 63180 489972 63232
rect 506296 63180 506348 63232
rect 547144 63180 547196 63232
rect 12348 63112 12400 63164
rect 62948 63112 63000 63164
rect 64144 63112 64196 63164
rect 83188 63112 83240 63164
rect 86868 63112 86920 63164
rect 123760 63112 123812 63164
rect 124128 63112 124180 63164
rect 154672 63112 154724 63164
rect 155868 63112 155920 63164
rect 180800 63112 180852 63164
rect 182088 63112 182140 63164
rect 202052 63112 202104 63164
rect 205548 63112 205600 63164
rect 221372 63112 221424 63164
rect 222108 63112 222160 63164
rect 234896 63112 234948 63164
rect 237288 63112 237340 63164
rect 247408 63112 247460 63164
rect 255964 63112 256016 63164
rect 261944 63112 261996 63164
rect 328552 63112 328604 63164
rect 329656 63112 329708 63164
rect 367192 63112 367244 63164
rect 368296 63112 368348 63164
rect 386512 63112 386564 63164
rect 387616 63112 387668 63164
rect 405832 63112 405884 63164
rect 406936 63112 406988 63164
rect 440608 63112 440660 63164
rect 441528 63112 441580 63164
rect 451280 63112 451332 63164
rect 467104 63112 467156 63164
rect 467656 63112 467708 63164
rect 502984 63112 503036 63164
rect 503444 63112 503496 63164
rect 544384 63112 544436 63164
rect 65524 63044 65576 63096
rect 89996 63044 90048 63096
rect 95148 63044 95200 63096
rect 131488 63044 131540 63096
rect 142068 63044 142120 63096
rect 169208 63044 169260 63096
rect 169668 63044 169720 63096
rect 192392 63044 192444 63096
rect 194416 63044 194468 63096
rect 211712 63044 211764 63096
rect 212448 63044 212500 63096
rect 227168 63044 227220 63096
rect 227628 63044 227680 63096
rect 239680 63044 239732 63096
rect 241428 63044 241480 63096
rect 250352 63044 250404 63096
rect 251088 63044 251140 63096
rect 258080 63044 258132 63096
rect 267648 63044 267700 63096
rect 271604 63044 271656 63096
rect 422300 63044 422352 63096
rect 436652 63044 436704 63096
rect 444472 63044 444524 63096
rect 464344 63044 464396 63096
rect 474464 63044 474516 63096
rect 490564 63044 490616 63096
rect 490840 63044 490892 63096
rect 532056 63044 532108 63096
rect 16488 62976 16540 63028
rect 66812 62976 66864 63028
rect 72424 62976 72476 63028
rect 78404 62976 78456 63028
rect 13728 62908 13780 62960
rect 64880 62908 64932 62960
rect 71688 62908 71740 62960
rect 81348 62976 81400 63028
rect 119896 62976 119948 63028
rect 119988 62976 120040 63028
rect 151820 62976 151872 63028
rect 153108 62976 153160 63028
rect 178868 62976 178920 63028
rect 179328 62976 179380 63028
rect 200120 62976 200172 63028
rect 206928 62976 206980 63028
rect 222292 62976 222344 63028
rect 224868 62976 224920 63028
rect 236828 62976 236880 63028
rect 238668 62976 238720 63028
rect 248420 62976 248472 63028
rect 257988 62976 258040 63028
rect 263876 62976 263928 63028
rect 311164 62976 311216 63028
rect 311808 62976 311860 63028
rect 318892 62976 318944 63028
rect 321008 62976 321060 63028
rect 330484 62976 330536 63028
rect 331128 62976 331180 63028
rect 349804 62976 349856 63028
rect 350448 62976 350500 63028
rect 369124 62976 369176 63028
rect 369768 62976 369820 63028
rect 388444 62976 388496 63028
rect 389088 62976 389140 63028
rect 407764 62976 407816 63028
rect 408408 62976 408460 63028
rect 421288 62976 421340 63028
rect 422208 62976 422260 63028
rect 427084 62976 427136 63028
rect 427728 62976 427780 63028
rect 437756 62976 437808 63028
rect 454684 62976 454736 63028
rect 463792 62976 463844 63028
rect 500316 62976 500368 63028
rect 500500 62976 500552 63028
rect 543004 62976 543056 63028
rect 6828 62840 6880 62892
rect 59084 62840 59136 62892
rect 62764 62840 62816 62892
rect 70676 62840 70728 62892
rect 73804 62840 73856 62892
rect 76472 62840 76524 62892
rect 76564 62840 76616 62892
rect 85120 62908 85172 62960
rect 88248 62908 88300 62960
rect 125692 62908 125744 62960
rect 129004 62908 129056 62960
rect 138296 62908 138348 62960
rect 143448 62908 143500 62960
rect 170128 62908 170180 62960
rect 171048 62908 171100 62960
rect 193312 62908 193364 62960
rect 194508 62908 194560 62960
rect 212632 62908 212684 62960
rect 213828 62908 213880 62960
rect 228088 62908 228140 62960
rect 230388 62908 230440 62960
rect 241612 62908 241664 62960
rect 242808 62908 242860 62960
rect 251272 62908 251324 62960
rect 267004 62908 267056 62960
rect 270592 62908 270644 62960
rect 423220 62908 423272 62960
rect 112168 62840 112220 62892
rect 113088 62840 113140 62892
rect 146024 62840 146076 62892
rect 150348 62840 150400 62892
rect 175924 62840 175976 62892
rect 177856 62840 177908 62892
rect 199108 62840 199160 62892
rect 202696 62840 202748 62892
rect 219440 62840 219492 62892
rect 220728 62840 220780 62892
rect 233884 62840 233936 62892
rect 234528 62840 234580 62892
rect 244556 62840 244608 62892
rect 245568 62840 245620 62892
rect 254216 62840 254268 62892
rect 256608 62840 256660 62892
rect 262864 62840 262916 62892
rect 327632 62840 327684 62892
rect 328368 62840 328420 62892
rect 346952 62840 347004 62892
rect 347688 62840 347740 62892
rect 366272 62840 366324 62892
rect 367008 62840 367060 62892
rect 385592 62840 385644 62892
rect 386328 62840 386380 62892
rect 404912 62840 404964 62892
rect 405648 62840 405700 62892
rect 416504 62840 416556 62892
rect 4068 62772 4120 62824
rect 57152 62772 57204 62824
rect 57888 62772 57940 62824
rect 100576 62772 100628 62824
rect 103428 62772 103480 62824
rect 137284 62772 137336 62824
rect 139308 62772 139360 62824
rect 167276 62772 167328 62824
rect 168288 62772 168340 62824
rect 190460 62772 190512 62824
rect 191748 62772 191800 62824
rect 209780 62772 209832 62824
rect 210976 62772 211028 62824
rect 226156 62772 226208 62824
rect 227536 62772 227588 62824
rect 238760 62772 238812 62824
rect 244096 62772 244148 62824
rect 253204 62772 253256 62824
rect 253848 62772 253900 62824
rect 260932 62772 260984 62824
rect 277216 62772 277268 62824
rect 280252 62772 280304 62824
rect 340144 62772 340196 62824
rect 340788 62772 340840 62824
rect 359464 62772 359516 62824
rect 360108 62772 360160 62824
rect 378784 62772 378836 62824
rect 379428 62772 379480 62824
rect 398104 62772 398156 62824
rect 398748 62772 398800 62824
rect 417424 62772 417476 62824
rect 418068 62772 418120 62824
rect 424232 62840 424284 62892
rect 424968 62840 425020 62892
rect 434812 62908 434864 62960
rect 465172 62908 465224 62960
rect 468668 62908 468720 62960
rect 487804 62908 487856 62960
rect 491852 62908 491904 62960
rect 535460 62908 535512 62960
rect 446312 62840 446364 62892
rect 464804 62840 464856 62892
rect 431224 62772 431276 62824
rect 442540 62772 442592 62824
rect 474004 62772 474056 62824
rect 492772 62840 492824 62892
rect 493968 62840 494020 62892
rect 497648 62840 497700 62892
rect 541624 62840 541676 62892
rect 497464 62772 497516 62824
rect 529204 62772 529256 62824
rect 529480 62772 529532 62824
rect 33048 62704 33100 62756
rect 80336 62704 80388 62756
rect 80704 62704 80756 62756
rect 90916 62704 90968 62756
rect 91744 62704 91796 62756
rect 108304 62704 108356 62756
rect 117228 62704 117280 62756
rect 148876 62704 148928 62756
rect 162768 62704 162820 62756
rect 186596 62704 186648 62756
rect 188988 62704 189040 62756
rect 207848 62704 207900 62756
rect 208308 62704 208360 62756
rect 223304 62704 223356 62756
rect 235816 62704 235868 62756
rect 245476 62704 245528 62756
rect 302516 62704 302568 62756
rect 303344 62704 303396 62756
rect 325700 62704 325752 62756
rect 331864 62704 331916 62756
rect 486056 62704 486108 62756
rect 525064 62704 525116 62756
rect 528560 62704 528612 62756
rect 545764 62704 545816 62756
rect 39948 62636 40000 62688
rect 86132 62636 86184 62688
rect 122748 62636 122800 62688
rect 153752 62636 153804 62688
rect 158628 62636 158680 62688
rect 182732 62636 182784 62688
rect 190368 62636 190420 62688
rect 208768 62636 208820 62688
rect 217968 62636 218020 62688
rect 231032 62636 231084 62688
rect 313096 62636 313148 62688
rect 313924 62636 313976 62688
rect 351736 62636 351788 62688
rect 352564 62636 352616 62688
rect 487988 62636 488040 62688
rect 526444 62636 526496 62688
rect 34428 62568 34480 62620
rect 81256 62568 81308 62620
rect 97264 62568 97316 62620
rect 106372 62568 106424 62620
rect 107016 62568 107068 62620
rect 122840 62568 122892 62620
rect 125508 62568 125560 62620
rect 155684 62568 155736 62620
rect 160008 62568 160060 62620
rect 183652 62568 183704 62620
rect 184848 62568 184900 62620
rect 203984 62568 204036 62620
rect 219348 62568 219400 62620
rect 232964 62568 233016 62620
rect 452200 62568 452252 62620
rect 453304 62568 453356 62620
rect 477316 62568 477368 62620
rect 515496 62568 515548 62620
rect 515956 62568 516008 62620
rect 517520 62568 517572 62620
rect 523684 62568 523736 62620
rect 551284 62568 551336 62620
rect 41328 62500 41380 62552
rect 87052 62500 87104 62552
rect 95884 62500 95936 62552
rect 111248 62500 111300 62552
rect 116584 62500 116636 62552
rect 143080 62500 143132 62552
rect 146944 62500 146996 62552
rect 158536 62500 158588 62552
rect 164148 62500 164200 62552
rect 187516 62500 187568 62552
rect 187608 62500 187660 62552
rect 206836 62500 206888 62552
rect 216588 62500 216640 62552
rect 230020 62500 230072 62552
rect 478328 62500 478380 62552
rect 479524 62500 479576 62552
rect 50988 62432 51040 62484
rect 94780 62432 94832 62484
rect 100116 62432 100168 62484
rect 109316 62432 109368 62484
rect 112444 62432 112496 62484
rect 128636 62432 128688 62484
rect 137284 62432 137336 62484
rect 149888 62432 149940 62484
rect 161388 62432 161440 62484
rect 184664 62432 184716 62484
rect 195888 62432 195940 62484
rect 213644 62432 213696 62484
rect 321836 62432 321888 62484
rect 322848 62432 322900 62484
rect 333428 62432 333480 62484
rect 334624 62432 334676 62484
rect 391388 62432 391440 62484
rect 392584 62432 392636 62484
rect 476396 62432 476448 62484
rect 513932 62500 513984 62552
rect 519820 62500 519872 62552
rect 534724 62500 534776 62552
rect 505376 62432 505428 62484
rect 540336 62432 540388 62484
rect 43444 62364 43496 62416
rect 79324 62364 79376 62416
rect 113824 62364 113876 62416
rect 126704 62364 126756 62416
rect 135904 62364 135956 62416
rect 146852 62364 146904 62416
rect 156604 62364 156656 62416
rect 164332 62364 164384 62416
rect 166908 62364 166960 62416
rect 189448 62364 189500 62416
rect 193128 62364 193180 62416
rect 210700 62364 210752 62416
rect 260748 62364 260800 62416
rect 266728 62364 266780 62416
rect 308312 62364 308364 62416
rect 309784 62364 309836 62416
rect 341156 62364 341208 62416
rect 342168 62364 342220 62416
rect 360476 62364 360528 62416
rect 361488 62364 361540 62416
rect 399116 62364 399168 62416
rect 400128 62364 400180 62416
rect 418436 62364 418488 62416
rect 419448 62364 419500 62416
rect 420368 62364 420420 62416
rect 421564 62364 421616 62416
rect 441620 62364 441672 62416
rect 442908 62364 442960 62416
rect 483112 62364 483164 62416
rect 515404 62364 515456 62416
rect 525616 62364 525668 62416
rect 540244 62364 540296 62416
rect 53104 62296 53156 62348
rect 93860 62296 93912 62348
rect 108304 62296 108356 62348
rect 117964 62296 118016 62348
rect 123484 62296 123536 62348
rect 135352 62296 135404 62348
rect 160744 62296 160796 62348
rect 173072 62296 173124 62348
rect 173808 62296 173860 62348
rect 195244 62296 195296 62348
rect 200028 62296 200080 62348
rect 216496 62296 216548 62348
rect 259368 62296 259420 62348
rect 264796 62296 264848 62348
rect 269028 62296 269080 62348
rect 273536 62296 273588 62348
rect 316040 62296 316092 62348
rect 317328 62296 317380 62348
rect 335360 62296 335412 62348
rect 336648 62296 336700 62348
rect 338212 62296 338264 62348
rect 339408 62296 339460 62348
rect 357532 62296 357584 62348
rect 358728 62296 358780 62348
rect 374000 62296 374052 62348
rect 375288 62296 375340 62348
rect 376852 62296 376904 62348
rect 378048 62296 378100 62348
rect 379796 62296 379848 62348
rect 381544 62296 381596 62348
rect 393320 62296 393372 62348
rect 394608 62296 394660 62348
rect 396172 62296 396224 62348
rect 397368 62296 397420 62348
rect 524696 62296 524748 62348
rect 531964 62296 532016 62348
rect 15108 62228 15160 62280
rect 65800 62228 65852 62280
rect 66904 62228 66956 62280
rect 96712 62228 96764 62280
rect 98644 62228 98696 62280
rect 114100 62228 114152 62280
rect 120724 62228 120776 62280
rect 132500 62228 132552 62280
rect 176568 62228 176620 62280
rect 197176 62228 197228 62280
rect 201408 62228 201460 62280
rect 217508 62228 217560 62280
rect 249708 62228 249760 62280
rect 257068 62228 257120 62280
rect 263508 62228 263560 62280
rect 268660 62228 268712 62280
rect 270408 62228 270460 62280
rect 274456 62228 274508 62280
rect 274548 62228 274600 62280
rect 277400 62228 277452 62280
rect 319904 62228 319956 62280
rect 320916 62228 320968 62280
rect 408776 62228 408828 62280
rect 410524 62228 410576 62280
rect 450268 62228 450320 62280
rect 451188 62228 451240 62280
rect 481180 62228 481232 62280
rect 485136 62228 485188 62280
rect 55864 62160 55916 62212
rect 84200 62160 84252 62212
rect 106924 62160 106976 62212
rect 115112 62160 115164 62212
rect 133144 62160 133196 62212
rect 141148 62160 141200 62212
rect 188344 62160 188396 62212
rect 204904 62160 204956 62212
rect 252376 62160 252428 62212
rect 260012 62160 260064 62212
rect 264888 62160 264940 62212
rect 269672 62160 269724 62212
rect 271788 62160 271840 62212
rect 275468 62160 275520 62212
rect 275928 62160 275980 62212
rect 278320 62160 278372 62212
rect 278688 62160 278740 62212
rect 281264 62160 281316 62212
rect 281448 62160 281500 62212
rect 283196 62160 283248 62212
rect 315028 62160 315080 62212
rect 318064 62160 318116 62212
rect 433892 62160 433944 62212
rect 439504 62160 439556 62212
rect 469588 62160 469640 62212
rect 472624 62160 472676 62212
rect 473452 62160 473504 62212
rect 476764 62160 476816 62212
rect 480260 62160 480312 62212
rect 483664 62160 483716 62212
rect 510160 62160 510212 62212
rect 511264 62160 511316 62212
rect 60004 62092 60056 62144
rect 61016 62092 61068 62144
rect 61384 62092 61436 62144
rect 75184 62092 75236 62144
rect 82268 62092 82320 62144
rect 88984 62092 89036 62144
rect 91928 62092 91980 62144
rect 100024 62092 100076 62144
rect 103520 62092 103572 62144
rect 113916 62092 113968 62144
rect 120908 62092 120960 62144
rect 134616 62092 134668 62144
rect 136364 62092 136416 62144
rect 137376 62092 137428 62144
rect 139216 62092 139268 62144
rect 202788 62092 202840 62144
rect 218428 62092 218480 62144
rect 252468 62092 252520 62144
rect 259000 62092 259052 62144
rect 260656 62092 260708 62144
rect 265808 62092 265860 62144
rect 267096 62092 267148 62144
rect 267740 62092 267792 62144
rect 269764 62092 269816 62144
rect 272524 62092 272576 62144
rect 277308 62092 277360 62144
rect 279332 62092 279384 62144
rect 280804 62092 280856 62144
rect 282184 62092 282236 62144
rect 282828 62092 282880 62144
rect 284116 62092 284168 62144
rect 285588 62092 285640 62144
rect 287060 62092 287112 62144
rect 288348 62092 288400 62144
rect 288992 62092 289044 62144
rect 289820 62092 289872 62144
rect 290924 62092 290976 62144
rect 292580 62092 292632 62144
rect 293776 62092 293828 62144
rect 297640 62092 297692 62144
rect 298192 62092 298244 62144
rect 298652 62092 298704 62144
rect 299388 62092 299440 62144
rect 301504 62092 301556 62144
rect 302424 62092 302476 62144
rect 304448 62092 304500 62144
rect 304908 62092 304960 62144
rect 305368 62092 305420 62144
rect 306288 62092 306340 62144
rect 306380 62092 306432 62144
rect 307668 62092 307720 62144
rect 309232 62092 309284 62144
rect 310336 62092 310388 62144
rect 312176 62092 312228 62144
rect 313188 62092 313240 62144
rect 314108 62092 314160 62144
rect 314568 62092 314620 62144
rect 317972 62092 318024 62144
rect 318708 62092 318760 62144
rect 320824 62092 320876 62144
rect 321468 62092 321520 62144
rect 323768 62092 323820 62144
rect 324228 62092 324280 62144
rect 324688 62092 324740 62144
rect 325608 62092 325660 62144
rect 331496 62092 331548 62144
rect 332324 62092 332376 62144
rect 337292 62092 337344 62144
rect 340236 62092 340288 62144
rect 343088 62092 343140 62144
rect 343548 62092 343600 62144
rect 344008 62092 344060 62144
rect 344928 62092 344980 62144
rect 345020 62092 345072 62144
rect 346216 62092 346268 62144
rect 347872 62092 347924 62144
rect 349068 62092 349120 62144
rect 350816 62092 350868 62144
rect 351828 62092 351880 62144
rect 352748 62092 352800 62144
rect 353208 62092 353260 62144
rect 354680 62092 354732 62144
rect 355876 62092 355928 62144
rect 356612 62092 356664 62144
rect 357348 62092 357400 62144
rect 362408 62092 362460 62144
rect 362868 62092 362920 62144
rect 363328 62092 363380 62144
rect 364248 62092 364300 62144
rect 364340 62092 364392 62144
rect 365628 62092 365680 62144
rect 370136 62092 370188 62144
rect 371148 62092 371200 62144
rect 372068 62092 372120 62144
rect 372528 62092 372580 62144
rect 375932 62092 375984 62144
rect 376668 62092 376720 62144
rect 381728 62092 381780 62144
rect 382188 62092 382240 62144
rect 382648 62092 382700 62144
rect 383568 62092 383620 62144
rect 383660 62092 383712 62144
rect 384856 62092 384908 62144
rect 389456 62092 389508 62144
rect 390284 62092 390336 62144
rect 395252 62092 395304 62144
rect 395988 62092 396040 62144
rect 401048 62092 401100 62144
rect 401508 62092 401560 62144
rect 401968 62092 402020 62144
rect 402888 62092 402940 62144
rect 402980 62092 403032 62144
rect 404176 62092 404228 62144
rect 410708 62092 410760 62144
rect 411168 62092 411220 62144
rect 412640 62092 412692 62144
rect 413836 62092 413888 62144
rect 414572 62092 414624 62144
rect 415308 62092 415360 62144
rect 415492 62092 415544 62144
rect 416688 62092 416740 62144
rect 425152 62092 425204 62144
rect 426348 62092 426400 62144
rect 428096 62092 428148 62144
rect 429108 62092 429160 62144
rect 430028 62092 430080 62144
rect 430488 62092 430540 62144
rect 430948 62092 431000 62144
rect 431868 62092 431920 62144
rect 431960 62092 432012 62144
rect 433156 62092 433208 62144
rect 436744 62092 436796 62144
rect 437388 62092 437440 62144
rect 443552 62092 443604 62144
rect 444288 62092 444340 62144
rect 446404 62092 446456 62144
rect 447048 62092 447100 62144
rect 447416 62092 447468 62144
rect 448244 62092 448296 62144
rect 449348 62092 449400 62144
rect 449808 62092 449860 62144
rect 453212 62092 453264 62144
rect 453948 62092 454000 62144
rect 456064 62092 456116 62144
rect 456708 62092 456760 62144
rect 459008 62092 459060 62144
rect 459468 62092 459520 62144
rect 459928 62092 459980 62144
rect 460848 62092 460900 62144
rect 460940 62092 460992 62144
rect 462136 62092 462188 62144
rect 465724 62092 465776 62144
rect 466368 62092 466420 62144
rect 466736 62092 466788 62144
rect 467748 62092 467800 62144
rect 472532 62092 472584 62144
rect 473268 62092 473320 62144
rect 475384 62092 475436 62144
rect 476028 62092 476080 62144
rect 479248 62092 479300 62144
rect 480168 62092 480220 62144
rect 485044 62092 485096 62144
rect 485688 62092 485740 62144
rect 488908 62092 488960 62144
rect 489828 62092 489880 62144
rect 495716 62092 495768 62144
rect 497556 62092 497608 62144
rect 498568 62092 498620 62144
rect 500224 62092 500276 62144
rect 501512 62092 501564 62144
rect 502248 62092 502300 62144
rect 502432 62092 502484 62144
rect 503628 62092 503680 62144
rect 504364 62092 504416 62144
rect 505008 62092 505060 62144
rect 507308 62092 507360 62144
rect 507768 62092 507820 62144
rect 508228 62092 508280 62144
rect 509148 62092 509200 62144
rect 511172 62092 511224 62144
rect 511908 62092 511960 62144
rect 512092 62092 512144 62144
rect 513196 62092 513248 62144
rect 514024 62092 514076 62144
rect 514668 62092 514720 62144
rect 515036 62092 515088 62144
rect 516048 62092 516100 62144
rect 516968 62092 517020 62144
rect 517428 62092 517480 62144
rect 517888 62092 517940 62144
rect 518808 62092 518860 62144
rect 518900 62092 518952 62144
rect 520188 62092 520240 62144
rect 520832 62092 520884 62144
rect 521568 62092 521620 62144
rect 526628 62092 526680 62144
rect 527088 62092 527140 62144
rect 527548 62092 527600 62144
rect 528468 62092 528520 62144
rect 36544 61956 36596 62008
rect 55220 61956 55272 62008
rect 91008 61956 91060 62008
rect 127624 61956 127676 62008
rect 151084 61956 151136 62008
rect 162400 61956 162452 62008
rect 29736 61888 29788 61940
rect 63868 61888 63920 61940
rect 84108 61888 84160 61940
rect 121828 61888 121880 61940
rect 141424 61888 141476 61940
rect 165344 61888 165396 61940
rect 35256 61820 35308 61872
rect 75460 61820 75512 61872
rect 79968 61820 80020 61872
rect 118976 61820 119028 61872
rect 151728 61820 151780 61872
rect 176936 61820 176988 61872
rect 52368 61752 52420 61804
rect 95792 61752 95844 61804
rect 97908 61752 97960 61804
rect 133420 61752 133472 61804
rect 147588 61752 147640 61804
rect 173992 61752 174044 61804
rect 18604 61684 18656 61736
rect 54300 61684 54352 61736
rect 55128 61684 55180 61736
rect 98552 61684 98604 61736
rect 140688 61684 140740 61736
rect 168196 61684 168248 61736
rect 48228 61616 48280 61668
rect 92848 61616 92900 61668
rect 95056 61616 95108 61668
rect 130568 61616 130620 61668
rect 22008 61548 22060 61600
rect 71596 61548 71648 61600
rect 77208 61548 77260 61600
rect 116032 61548 116084 61600
rect 133236 61548 133288 61600
rect 161480 61548 161532 61600
rect 17868 61480 17920 61532
rect 67732 61480 67784 61532
rect 70308 61480 70360 61532
rect 110236 61480 110288 61532
rect 131028 61480 131080 61532
rect 160468 61480 160520 61532
rect 165528 61480 165580 61532
rect 188528 61480 188580 61532
rect 517520 61480 517572 61532
rect 564532 61480 564584 61532
rect 4896 61412 4948 61464
rect 56140 61412 56192 61464
rect 73068 61412 73120 61464
rect 113180 61412 113232 61464
rect 126888 61412 126940 61464
rect 156512 61412 156564 61464
rect 162124 61412 162176 61464
rect 185584 61412 185636 61464
rect 513104 61412 513156 61464
rect 561680 61412 561732 61464
rect 8208 61344 8260 61396
rect 59912 61344 59964 61396
rect 66168 61344 66220 61396
rect 107384 61344 107436 61396
rect 111708 61344 111760 61396
rect 144644 61344 144696 61396
rect 144736 61344 144788 61396
rect 171140 61344 171192 61396
rect 173164 61344 173216 61396
rect 194324 61344 194376 61396
rect 521752 61344 521804 61396
rect 572812 61344 572864 61396
rect 130384 61276 130436 61328
rect 157616 61276 157668 61328
rect 155224 61208 155276 61260
rect 163412 61208 163464 61260
rect 533344 60664 533396 60716
rect 580172 60664 580224 60716
rect 2780 58896 2832 58948
rect 4804 58896 4856 58948
rect 556804 46860 556856 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 33784 45500 33836 45552
rect 3516 33056 3568 33108
rect 29644 33056 29696 33108
rect 558184 33056 558236 33108
rect 580172 33056 580224 33108
rect 511264 32376 511316 32428
rect 557540 32376 557592 32428
rect 560944 20612 560996 20664
rect 579988 20612 580040 20664
rect 292580 11704 292632 11756
rect 293684 11704 293736 11756
rect 479524 8916 479576 8968
rect 519544 8916 519596 8968
rect 520188 8916 520240 8968
rect 569132 8916 569184 8968
rect 3424 6808 3476 6860
rect 35164 6808 35216 6860
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 86776 6196 86828 6248
rect 124772 6196 124824 6248
rect 129372 6196 129424 6248
rect 159548 6196 159600 6248
rect 58440 6128 58492 6180
rect 101588 6128 101640 6180
rect 101036 6060 101088 6112
rect 134616 6128 134668 6180
rect 169760 6128 169812 6180
rect 191380 6128 191432 6180
rect 473268 6128 473320 6180
rect 512460 6128 512512 6180
rect 472624 5448 472676 5500
rect 508872 5448 508924 5500
rect 485136 5380 485188 5432
rect 523040 5380 523092 5432
rect 410524 5312 410576 5364
rect 434444 5312 434496 5364
rect 454684 5312 454736 5364
rect 469864 5312 469916 5364
rect 476028 5312 476080 5364
rect 515956 5312 516008 5364
rect 404176 5244 404228 5296
rect 427268 5244 427320 5296
rect 433156 5244 433208 5296
rect 462780 5244 462832 5296
rect 484308 5244 484360 5296
rect 526628 5244 526680 5296
rect 383568 5176 383620 5228
rect 402520 5176 402572 5228
rect 406936 5176 406988 5228
rect 430856 5176 430908 5228
rect 447048 5176 447100 5228
rect 480536 5176 480588 5228
rect 497556 5176 497608 5228
rect 540796 5176 540848 5228
rect 386328 5108 386380 5160
rect 406016 5108 406068 5160
rect 412548 5108 412600 5160
rect 437940 5108 437992 5160
rect 453304 5108 453356 5160
rect 487620 5108 487672 5160
rect 493968 5108 494020 5160
rect 537208 5108 537260 5160
rect 389088 5040 389140 5092
rect 409604 5040 409656 5092
rect 415308 5040 415360 5092
rect 441436 5040 441488 5092
rect 449808 5040 449860 5092
rect 484032 5040 484084 5092
rect 487068 5040 487120 5092
rect 530124 5040 530176 5092
rect 392584 4972 392636 5024
rect 413100 4972 413152 5024
rect 418068 4972 418120 5024
rect 445024 4972 445076 5024
rect 455328 4972 455380 5024
rect 491116 4972 491168 5024
rect 500224 4972 500276 5024
rect 544292 4972 544344 5024
rect 394516 4904 394568 4956
rect 416688 4904 416740 4956
rect 421564 4904 421616 4956
rect 448612 4904 448664 4956
rect 458088 4904 458140 4956
rect 494704 4904 494756 4956
rect 505008 4904 505060 4956
rect 551468 4904 551520 4956
rect 62028 4836 62080 4888
rect 104440 4836 104492 4888
rect 128360 4836 128412 4888
rect 142160 4836 142212 4888
rect 397276 4836 397328 4888
rect 420184 4836 420236 4888
rect 429016 4836 429068 4888
rect 459192 4836 459244 4888
rect 462136 4836 462188 4888
rect 498200 4836 498252 4888
rect 502248 4836 502300 4888
rect 547880 4836 547932 4888
rect 30104 4768 30156 4820
rect 72424 4768 72476 4820
rect 139400 4768 139452 4820
rect 166264 4768 166316 4820
rect 381544 4768 381596 4820
rect 398932 4768 398984 4820
rect 400036 4768 400088 4820
rect 423772 4768 423824 4820
rect 426256 4768 426308 4820
rect 455696 4768 455748 4820
rect 467748 4768 467800 4820
rect 505376 4768 505428 4820
rect 507768 4768 507820 4820
rect 554964 4768 555016 4820
rect 446404 4360 446456 4412
rect 452108 4360 452160 4412
rect 442908 4156 442960 4208
rect 45468 4088 45520 4140
rect 80704 4088 80756 4140
rect 123392 4088 123444 4140
rect 161296 4088 161348 4140
rect 162124 4088 162176 4140
rect 322848 4088 322900 4140
rect 328000 4088 328052 4140
rect 342168 4088 342220 4140
rect 351644 4088 351696 4140
rect 355876 4088 355928 4140
rect 368204 4088 368256 4140
rect 373908 4088 373960 4140
rect 390652 4088 390704 4140
rect 397368 4088 397420 4140
rect 418988 4088 419040 4140
rect 419448 4088 419500 4140
rect 446220 4088 446272 4140
rect 500316 4156 500368 4208
rect 501788 4156 501840 4208
rect 529204 4156 529256 4208
rect 533712 4156 533764 4208
rect 451188 4088 451240 4140
rect 485228 4088 485280 4140
rect 487804 4088 487856 4140
rect 507676 4088 507728 4140
rect 511908 4088 511960 4140
rect 559748 4088 559800 4140
rect 31300 4020 31352 4072
rect 43444 4020 43496 4072
rect 53748 4020 53800 4072
rect 90272 4020 90324 4072
rect 96252 4020 96304 4072
rect 120724 4020 120776 4072
rect 344928 4020 344980 4072
rect 355232 4020 355284 4072
rect 358728 4020 358780 4072
rect 371700 4020 371752 4072
rect 375196 4020 375248 4072
rect 393044 4020 393096 4072
rect 394608 4020 394660 4072
rect 415492 4020 415544 4072
rect 422208 4020 422260 4072
rect 449808 4020 449860 4072
rect 456708 4020 456760 4072
rect 492312 4020 492364 4072
rect 509148 4020 509200 4072
rect 556160 4020 556212 4072
rect 41880 3952 41932 4004
rect 79324 3952 79376 4004
rect 89168 3952 89220 4004
rect 113824 3952 113876 4004
rect 128176 3952 128228 4004
rect 146944 3952 146996 4004
rect 334624 3952 334676 4004
rect 342168 3952 342220 4004
rect 343548 3952 343600 4004
rect 354036 3952 354088 4004
rect 355968 3952 356020 4004
rect 369400 3952 369452 4004
rect 372528 3952 372580 4004
rect 389456 3952 389508 4004
rect 390284 3952 390336 4004
rect 410800 3952 410852 4004
rect 413928 3952 413980 4004
rect 439504 3952 439556 4004
rect 38384 3884 38436 3936
rect 77392 3884 77444 3936
rect 99840 3884 99892 3936
rect 12256 3816 12308 3868
rect 29736 3816 29788 3868
rect 34796 3816 34848 3868
rect 75184 3816 75236 3868
rect 78588 3816 78640 3868
rect 20536 3748 20588 3800
rect 62764 3748 62816 3800
rect 1676 3680 1728 3732
rect 36544 3680 36596 3732
rect 50160 3680 50212 3732
rect 50988 3680 51040 3732
rect 51356 3680 51408 3732
rect 52368 3680 52420 3732
rect 76564 3748 76616 3800
rect 88984 3680 89036 3732
rect 105544 3748 105596 3800
rect 108120 3816 108172 3868
rect 128360 3884 128412 3936
rect 349068 3884 349120 3936
rect 359924 3884 359976 3936
rect 362868 3884 362920 3936
rect 377680 3884 377732 3936
rect 379428 3884 379480 3936
rect 397736 3884 397788 3936
rect 398748 3884 398800 3936
rect 421380 3884 421432 3936
rect 426348 3884 426400 3936
rect 453948 3952 454000 4004
rect 488816 3952 488868 4004
rect 513196 3952 513248 4004
rect 560852 3952 560904 4004
rect 465172 3884 465224 3936
rect 109316 3816 109368 3868
rect 116584 3816 116636 3868
rect 117596 3816 117648 3868
rect 137284 3816 137336 3868
rect 314568 3816 314620 3868
rect 318524 3816 318576 3868
rect 336556 3816 336608 3868
rect 346216 3816 346268 3868
rect 356336 3816 356388 3868
rect 360108 3816 360160 3868
rect 374092 3816 374144 3868
rect 380808 3816 380860 3868
rect 400036 3816 400088 3868
rect 400128 3816 400180 3868
rect 422576 3816 422628 3868
rect 424968 3816 425020 3868
rect 453304 3816 453356 3868
rect 460388 3816 460440 3868
rect 460848 3816 460900 3868
rect 497096 3884 497148 3936
rect 514668 3884 514720 3936
rect 563244 3884 563296 3936
rect 108304 3748 108356 3800
rect 114008 3748 114060 3800
rect 135904 3748 135956 3800
rect 335268 3748 335320 3800
rect 343364 3748 343416 3800
rect 350356 3748 350408 3800
rect 362316 3748 362368 3800
rect 367008 3748 367060 3800
rect 382372 3748 382424 3800
rect 384856 3748 384908 3800
rect 403624 3748 403676 3800
rect 404268 3748 404320 3800
rect 428464 3748 428516 3800
rect 430488 3748 430540 3800
rect 454500 3748 454552 3800
rect 495900 3816 495952 3868
rect 497464 3816 497516 3868
rect 502892 3816 502944 3868
rect 516048 3816 516100 3868
rect 564440 3816 564492 3868
rect 100116 3680 100168 3732
rect 103336 3680 103388 3732
rect 129004 3680 129056 3732
rect 132960 3680 133012 3732
rect 151084 3680 151136 3732
rect 320916 3680 320968 3732
rect 325516 3680 325568 3732
rect 325608 3680 325660 3732
rect 331588 3680 331640 3732
rect 332324 3680 332376 3732
rect 339868 3680 339920 3732
rect 340788 3680 340840 3732
rect 350448 3680 350500 3732
rect 353208 3680 353260 3732
rect 365812 3680 365864 3732
rect 368388 3680 368440 3732
rect 384764 3680 384816 3732
rect 387616 3680 387668 3732
rect 407212 3680 407264 3732
rect 413836 3680 413888 3732
rect 439136 3680 439188 3732
rect 440148 3680 440200 3732
rect 572 3544 624 3596
rect 18604 3612 18656 3664
rect 8760 3544 8812 3596
rect 2872 3476 2924 3528
rect 4896 3476 4948 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 15936 3544 15988 3596
rect 16488 3544 16540 3596
rect 17040 3544 17092 3596
rect 17868 3544 17920 3596
rect 18236 3544 18288 3596
rect 19432 3544 19484 3596
rect 20628 3544 20680 3596
rect 24216 3544 24268 3596
rect 24768 3544 24820 3596
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 68744 3612 68796 3664
rect 73804 3612 73856 3664
rect 75000 3612 75052 3664
rect 106924 3612 106976 3664
rect 110512 3612 110564 3664
rect 134524 3612 134576 3664
rect 65524 3544 65576 3596
rect 66168 3544 66220 3596
rect 69112 3544 69164 3596
rect 70308 3544 70360 3596
rect 72608 3544 72660 3596
rect 73068 3544 73120 3596
rect 76196 3544 76248 3596
rect 77208 3544 77260 3596
rect 80888 3544 80940 3596
rect 81348 3544 81400 3596
rect 82084 3544 82136 3596
rect 113916 3544 113968 3596
rect 115204 3544 115256 3596
rect 115848 3544 115900 3596
rect 116400 3544 116452 3596
rect 117228 3544 117280 3596
rect 118792 3544 118844 3596
rect 119804 3544 119856 3596
rect 122288 3544 122340 3596
rect 122748 3544 122800 3596
rect 124680 3544 124732 3596
rect 125508 3544 125560 3596
rect 125876 3544 125928 3596
rect 126888 3544 126940 3596
rect 126980 3544 127032 3596
rect 130384 3544 130436 3596
rect 130568 3544 130620 3596
rect 131028 3544 131080 3596
rect 134156 3544 134208 3596
rect 155224 3544 155276 3596
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 64328 3476 64380 3528
rect 5264 3408 5316 3460
rect 58072 3408 58124 3460
rect 60832 3408 60884 3460
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 102232 3476 102284 3528
rect 103428 3476 103480 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 133144 3476 133196 3528
rect 97264 3408 97316 3460
rect 104532 3408 104584 3460
rect 137376 3476 137428 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 156604 3612 156656 3664
rect 171968 3612 172020 3664
rect 173164 3612 173216 3664
rect 324228 3612 324280 3664
rect 330392 3612 330444 3664
rect 331128 3612 331180 3664
rect 338672 3612 338724 3664
rect 339408 3612 339460 3664
rect 348056 3612 348108 3664
rect 348976 3612 349028 3664
rect 361120 3612 361172 3664
rect 361396 3612 361448 3664
rect 376484 3612 376536 3664
rect 382188 3612 382240 3664
rect 401324 3612 401376 3664
rect 402888 3612 402940 3664
rect 426164 3612 426216 3664
rect 427728 3612 427780 3664
rect 456892 3612 456944 3664
rect 459468 3612 459520 3664
rect 499396 3748 499448 3800
rect 518808 3748 518860 3800
rect 568028 3748 568080 3800
rect 462412 3612 462464 3664
rect 466368 3680 466420 3732
rect 476764 3680 476816 3732
rect 513564 3680 513616 3732
rect 517428 3680 517480 3732
rect 566832 3680 566884 3732
rect 300768 3544 300820 3596
rect 301964 3544 302016 3596
rect 303528 3544 303580 3596
rect 305552 3544 305604 3596
rect 310428 3544 310480 3596
rect 313832 3544 313884 3596
rect 317328 3544 317380 3596
rect 320916 3544 320968 3596
rect 336648 3544 336700 3596
rect 344560 3544 344612 3596
rect 345756 3544 345808 3596
rect 346308 3544 346360 3596
rect 357532 3544 357584 3596
rect 358636 3544 358688 3596
rect 372896 3544 372948 3596
rect 377956 3544 378008 3596
rect 396540 3544 396592 3596
rect 405648 3544 405700 3596
rect 429660 3544 429712 3596
rect 433248 3544 433300 3596
rect 463976 3544 464028 3596
rect 467104 3544 467156 3596
rect 467564 3544 467616 3596
rect 502984 3612 503036 3664
rect 506480 3612 506532 3664
rect 521568 3612 521620 3664
rect 571524 3612 571576 3664
rect 472256 3544 472308 3596
rect 135260 3408 135312 3460
rect 155408 3476 155460 3528
rect 155868 3476 155920 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 164884 3476 164936 3528
rect 165528 3476 165580 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 167184 3476 167236 3528
rect 168288 3476 168340 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 189724 3476 189776 3528
rect 190368 3476 190420 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 197912 3476 197964 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 200304 3476 200356 3528
rect 201408 3476 201460 3528
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 207388 3476 207440 3528
rect 208308 3476 208360 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 209780 3476 209832 3528
rect 211068 3476 211120 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 218060 3476 218112 3528
rect 219164 3476 219216 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 225144 3476 225196 3528
rect 226248 3476 226300 3528
rect 226340 3476 226392 3528
rect 227444 3476 227496 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235724 3476 235776 3528
rect 239312 3476 239364 3528
rect 240784 3476 240836 3528
rect 241704 3476 241756 3528
rect 242808 3476 242860 3528
rect 242900 3476 242952 3528
rect 244188 3476 244240 3528
rect 246396 3476 246448 3528
rect 246948 3476 247000 3528
rect 247592 3476 247644 3528
rect 248328 3476 248380 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 251180 3476 251232 3528
rect 252468 3476 252520 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 259460 3476 259512 3528
rect 260564 3476 260616 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 265348 3476 265400 3528
rect 267004 3476 267056 3528
rect 267740 3476 267792 3528
rect 269764 3476 269816 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 274824 3476 274876 3528
rect 275928 3476 275980 3528
rect 276020 3476 276072 3528
rect 277308 3476 277360 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 281908 3476 281960 3528
rect 282828 3476 282880 3528
rect 283104 3476 283156 3528
rect 285128 3476 285180 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 291384 3476 291436 3528
rect 291844 3476 291896 3528
rect 303344 3476 303396 3528
rect 304356 3476 304408 3528
rect 307668 3476 307720 3528
rect 309048 3476 309100 3528
rect 309784 3476 309836 3528
rect 311440 3476 311492 3528
rect 311808 3476 311860 3528
rect 315028 3476 315080 3528
rect 318064 3476 318116 3528
rect 319720 3476 319772 3528
rect 331864 3476 331916 3528
rect 332692 3476 332744 3528
rect 339316 3476 339368 3528
rect 349252 3476 349304 3528
rect 352564 3476 352616 3528
rect 364616 3476 364668 3528
rect 365536 3476 365588 3528
rect 381176 3476 381228 3528
rect 384948 3476 385000 3528
rect 404820 3476 404872 3528
rect 407028 3476 407080 3528
rect 432052 3476 432104 3528
rect 438768 3476 438820 3528
rect 471060 3476 471112 3528
rect 471888 3476 471940 3528
rect 511264 3544 511316 3596
rect 514024 3544 514076 3596
rect 517152 3544 517204 3596
rect 525064 3544 525116 3596
rect 529020 3544 529072 3596
rect 532056 3544 532108 3596
rect 534908 3544 534960 3596
rect 573916 3544 573968 3596
rect 474004 3476 474056 3528
rect 475752 3476 475804 3528
rect 480168 3476 480220 3528
rect 520740 3476 520792 3528
rect 527088 3476 527140 3528
rect 578608 3476 578660 3528
rect 141240 3408 141292 3460
rect 142068 3408 142120 3460
rect 142436 3408 142488 3460
rect 143448 3408 143500 3460
rect 143540 3408 143592 3460
rect 144644 3408 144696 3460
rect 147128 3408 147180 3460
rect 147588 3408 147640 3460
rect 148324 3408 148376 3460
rect 148968 3408 149020 3460
rect 149520 3408 149572 3460
rect 150348 3408 150400 3460
rect 150624 3408 150676 3460
rect 151728 3408 151780 3460
rect 240508 3408 240560 3460
rect 241428 3408 241480 3460
rect 248788 3408 248840 3460
rect 249708 3408 249760 3460
rect 254676 3408 254728 3460
rect 255964 3408 256016 3460
rect 266544 3408 266596 3460
rect 267648 3408 267700 3460
rect 286600 3408 286652 3460
rect 287980 3408 288032 3460
rect 304908 3408 304960 3460
rect 306748 3408 306800 3460
rect 307576 3408 307628 3460
rect 310244 3408 310296 3460
rect 322756 3408 322808 3460
rect 329196 3408 329248 3460
rect 332508 3408 332560 3460
rect 340972 3408 341024 3460
rect 342076 3408 342128 3460
rect 352840 3408 352892 3460
rect 357348 3408 357400 3460
rect 370596 3408 370648 3460
rect 371056 3408 371108 3460
rect 388260 3408 388312 3460
rect 390468 3408 390520 3460
rect 411904 3408 411956 3460
rect 419356 3408 419408 3460
rect 447416 3408 447468 3460
rect 448244 3408 448296 3460
rect 481732 3408 481784 3460
rect 485688 3408 485740 3460
rect 527824 3408 527876 3460
rect 528468 3408 528520 3460
rect 581000 3408 581052 3460
rect 25320 3340 25372 3392
rect 26148 3340 26200 3392
rect 27712 3340 27764 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 43076 3340 43128 3392
rect 77944 3340 77996 3392
rect 83280 3340 83332 3392
rect 84108 3340 84160 3392
rect 85672 3340 85724 3392
rect 86868 3340 86920 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 107016 3340 107068 3392
rect 121092 3340 121144 3392
rect 138664 3340 138716 3392
rect 145932 3340 145984 3392
rect 160744 3340 160796 3392
rect 313924 3340 313976 3392
rect 317328 3340 317380 3392
rect 351828 3340 351880 3392
rect 363512 3340 363564 3392
rect 369768 3340 369820 3392
rect 385960 3340 386012 3392
rect 387708 3340 387760 3392
rect 408408 3340 408460 3392
rect 409788 3340 409840 3392
rect 435548 3340 435600 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 473452 3340 473504 3392
rect 28908 3272 28960 3324
rect 35992 3204 36044 3256
rect 60004 3272 60056 3324
rect 70308 3272 70360 3324
rect 26516 3136 26568 3188
rect 35256 3136 35308 3188
rect 37188 3136 37240 3188
rect 48964 3136 49016 3188
rect 53104 3136 53156 3188
rect 55864 3068 55916 3120
rect 61384 3204 61436 3256
rect 64144 3204 64196 3256
rect 66720 3204 66772 3256
rect 95884 3272 95936 3324
rect 123484 3272 123536 3324
rect 124128 3272 124180 3324
rect 131764 3272 131816 3324
rect 133236 3272 133288 3324
rect 138848 3272 138900 3324
rect 139308 3272 139360 3324
rect 163688 3272 163740 3324
rect 164148 3272 164200 3324
rect 184940 3272 184992 3324
rect 188344 3272 188396 3324
rect 229836 3272 229888 3324
rect 230388 3272 230440 3324
rect 238116 3272 238168 3324
rect 238668 3272 238720 3324
rect 257068 3272 257120 3324
rect 257988 3272 258040 3324
rect 261760 3272 261812 3324
rect 267096 3272 267148 3324
rect 272432 3272 272484 3324
rect 276388 3272 276440 3324
rect 279516 3272 279568 3324
rect 280804 3272 280856 3324
rect 306288 3272 306340 3324
rect 307944 3272 307996 3324
rect 321008 3272 321060 3324
rect 324412 3272 324464 3324
rect 328368 3272 328420 3324
rect 335084 3272 335136 3324
rect 347688 3272 347740 3324
rect 358728 3272 358780 3324
rect 361488 3272 361540 3324
rect 375288 3272 375340 3324
rect 92756 3204 92808 3256
rect 93768 3204 93820 3256
rect 100024 3204 100076 3256
rect 136456 3204 136508 3256
rect 141424 3204 141476 3256
rect 318708 3204 318760 3256
rect 323308 3204 323360 3256
rect 354588 3204 354640 3256
rect 367008 3204 367060 3256
rect 375196 3204 375248 3256
rect 391848 3272 391900 3324
rect 393228 3272 393280 3324
rect 414296 3272 414348 3324
rect 416596 3272 416648 3324
rect 442632 3272 442684 3324
rect 444288 3272 444340 3324
rect 376668 3204 376720 3256
rect 394240 3204 394292 3256
rect 411168 3204 411220 3256
rect 436744 3204 436796 3256
rect 448428 3272 448480 3324
rect 482836 3340 482888 3392
rect 495348 3340 495400 3392
rect 539600 3340 539652 3392
rect 541624 3340 541676 3392
rect 543188 3340 543240 3392
rect 544384 3340 544436 3392
rect 482284 3272 482336 3324
rect 500592 3272 500644 3324
rect 504180 3272 504232 3324
rect 508504 3272 508556 3324
rect 510068 3272 510120 3324
rect 543004 3272 543056 3324
rect 546684 3272 546736 3324
rect 577412 3340 577464 3392
rect 550272 3272 550324 3324
rect 551284 3272 551336 3324
rect 575112 3272 575164 3324
rect 84844 3136 84896 3188
rect 91560 3136 91612 3188
rect 112444 3136 112496 3188
rect 193220 3136 193272 3188
rect 194324 3136 194376 3188
rect 216864 3136 216916 3188
rect 217968 3136 218020 3188
rect 310336 3136 310388 3188
rect 312636 3136 312688 3188
rect 317236 3136 317288 3188
rect 322112 3136 322164 3188
rect 329656 3136 329708 3188
rect 336280 3136 336332 3188
rect 378048 3136 378100 3188
rect 395344 3136 395396 3188
rect 408316 3136 408368 3188
rect 433248 3136 433300 3188
rect 436008 3136 436060 3188
rect 476948 3204 477000 3256
rect 489828 3204 489880 3256
rect 532516 3204 532568 3256
rect 533436 3204 533488 3256
rect 538404 3204 538456 3256
rect 467472 3136 467524 3188
rect 467564 3136 467616 3188
rect 486424 3136 486476 3188
rect 503628 3136 503680 3188
rect 63224 3068 63276 3120
rect 87604 3068 87656 3120
rect 168380 3068 168432 3120
rect 169760 3068 169812 3120
rect 221556 3068 221608 3120
rect 222108 3068 222160 3120
rect 313188 3068 313240 3120
rect 316224 3068 316276 3120
rect 340236 3068 340288 3120
rect 346952 3068 347004 3120
rect 371148 3068 371200 3120
rect 387156 3068 387208 3120
rect 401508 3068 401560 3120
rect 424968 3068 425020 3120
rect 437388 3068 437440 3120
rect 468668 3068 468720 3120
rect 478144 3068 478196 3120
rect 483664 3068 483716 3120
rect 522856 3136 522908 3188
rect 540336 3136 540388 3188
rect 521844 3068 521896 3120
rect 526444 3068 526496 3120
rect 531320 3068 531372 3120
rect 531964 3068 532016 3120
rect 576308 3204 576360 3256
rect 44272 3000 44324 3052
rect 65432 3000 65484 3052
rect 67916 3000 67968 3052
rect 46664 2932 46716 2984
rect 56048 2932 56100 2984
rect 73804 3000 73856 3052
rect 98552 3000 98604 3052
rect 151820 3000 151872 3052
rect 152924 3000 152976 3052
rect 196808 3000 196860 3052
rect 197268 3000 197320 3052
rect 321468 3000 321520 3052
rect 326804 3000 326856 3052
rect 329748 3000 329800 3052
rect 337476 3000 337528 3052
rect 368296 3000 368348 3052
rect 383568 3000 383620 3052
rect 395988 3000 396040 3052
rect 417884 3000 417936 3052
rect 431224 3000 431276 3052
rect 443828 3000 443880 3052
rect 449164 3000 449216 3052
rect 52552 2864 52604 2916
rect 66904 2864 66956 2916
rect 91744 2932 91796 2984
rect 284300 2932 284352 2984
rect 286048 2932 286100 2984
rect 326988 2932 327040 2984
rect 333888 2932 333940 2984
rect 365628 2932 365680 2984
rect 379980 2932 380032 2984
rect 436836 2932 436888 2984
rect 450912 2932 450964 2984
rect 474556 3000 474608 3052
rect 490564 3000 490616 3052
rect 514760 3000 514812 3052
rect 515496 3000 515548 3052
rect 518348 3000 518400 3052
rect 525432 3000 525484 3052
rect 534724 3000 534776 3052
rect 570328 3136 570380 3188
rect 545764 3068 545816 3120
rect 582196 3068 582248 3120
rect 552664 3000 552716 3052
rect 583392 3000 583444 3052
rect 479340 2932 479392 2984
rect 482928 2932 482980 2984
rect 524236 2932 524288 2984
rect 537484 2932 537536 2984
rect 541992 2932 542044 2984
rect 75276 2864 75328 2916
rect 84476 2864 84528 2916
rect 93952 2864 94004 2916
rect 95056 2864 95108 2916
rect 287796 2864 287848 2916
rect 288348 2864 288400 2916
rect 364248 2864 364300 2916
rect 378876 2864 378928 2916
rect 431868 2864 431920 2916
rect 461584 2864 461636 2916
rect 464344 2864 464396 2916
rect 471244 2864 471296 2916
rect 493508 2864 493560 2916
rect 515404 2864 515456 2916
rect 540244 2864 540296 2916
rect 548524 2932 548576 2984
rect 557356 2932 557408 2984
rect 549076 2864 549128 2916
rect 59636 2796 59688 2848
rect 137652 2796 137704 2848
rect 139400 2796 139452 2848
rect 429108 2796 429160 2848
rect 458088 2796 458140 2848
rect 468484 2796 468536 2848
rect 489920 2796 489972 2848
rect 538864 2796 538916 2848
rect 545488 2796 545540 2848
rect 547144 2796 547196 2848
rect 553768 2796 553820 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 105464 700534 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 166264 700528 166316 700534
rect 166264 700470 166316 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 166276 642462 166304 700470
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 235184 700534 235212 703520
rect 260748 700868 260800 700874
rect 260748 700810 260800 700816
rect 248328 700596 248380 700602
rect 248328 700538 248380 700544
rect 235172 700528 235224 700534
rect 235172 700470 235224 700476
rect 242164 700528 242216 700534
rect 242164 700470 242216 700476
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 171060 642530 171088 699654
rect 235908 696992 235960 696998
rect 235908 696934 235960 696940
rect 231768 670812 231820 670818
rect 231768 670754 231820 670760
rect 231780 644474 231808 670754
rect 231688 644446 231808 644474
rect 222936 643136 222988 643142
rect 222936 643078 222988 643084
rect 171048 642524 171100 642530
rect 171048 642466 171100 642472
rect 166264 642456 166316 642462
rect 166264 642398 166316 642404
rect 32404 641708 32456 641714
rect 32404 641650 32456 641656
rect 14464 641096 14516 641102
rect 14464 641038 14516 641044
rect 4802 640792 4858 640801
rect 4802 640727 4858 640736
rect 3516 638648 3568 638654
rect 3516 638590 3568 638596
rect 3422 638208 3478 638217
rect 3422 638143 3478 638152
rect 3332 632324 3384 632330
rect 3332 632266 3384 632272
rect 3344 632097 3372 632266
rect 3330 632088 3386 632097
rect 3330 632023 3386 632032
rect 3056 607164 3108 607170
rect 3056 607106 3108 607112
rect 3068 606121 3096 607106
rect 3054 606112 3110 606121
rect 3054 606047 3110 606056
rect 3332 580984 3384 580990
rect 3332 580926 3384 580932
rect 3344 580009 3372 580926
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3332 567180 3384 567186
rect 3332 567122 3384 567128
rect 3344 566953 3372 567122
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3332 554736 3384 554742
rect 3332 554678 3384 554684
rect 3344 553897 3372 554678
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3332 528556 3384 528562
rect 3332 528498 3384 528504
rect 3344 527921 3372 528498
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3148 516112 3200 516118
rect 3148 516054 3200 516060
rect 3160 514865 3188 516054
rect 3146 514856 3202 514865
rect 3146 514791 3202 514800
rect 2964 502308 3016 502314
rect 2964 502250 3016 502256
rect 2976 501809 3004 502250
rect 2962 501800 3018 501809
rect 2962 501735 3018 501744
rect 3240 476060 3292 476066
rect 3240 476002 3292 476008
rect 3252 475697 3280 476002
rect 3238 475688 3294 475697
rect 3238 475623 3294 475632
rect 3056 463684 3108 463690
rect 3056 463626 3108 463632
rect 3068 462641 3096 463626
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3332 372564 3384 372570
rect 3332 372506 3384 372512
rect 3344 371385 3372 372506
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 58948 2832 58954
rect 2780 58890 2832 58896
rect 2792 58585 2820 58890
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 3436 19417 3464 638143
rect 3528 201929 3556 638590
rect 3608 619608 3660 619614
rect 3608 619550 3660 619556
rect 3620 619177 3648 619550
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 188896 3568 188902
rect 3514 188864 3516 188873
rect 3568 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 4068 62824 4120 62830
rect 4068 62766 4120 62772
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 572 3596 624 3602
rect 572 3538 624 3544
rect 584 480 612 3538
rect 1688 480 1716 3674
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 480 2912 3470
rect 4080 480 4108 62766
rect 4816 58954 4844 640727
rect 7656 640008 7708 640014
rect 7656 639950 7708 639956
rect 7564 637764 7616 637770
rect 7564 637706 7616 637712
rect 7576 188902 7604 637706
rect 7668 632330 7696 639950
rect 11796 639940 11848 639946
rect 11796 639882 11848 639888
rect 11702 637664 11758 637673
rect 11702 637599 11758 637608
rect 7656 632324 7708 632330
rect 7656 632266 7708 632272
rect 7564 188896 7616 188902
rect 7564 188838 7616 188844
rect 11716 85542 11744 637599
rect 11808 580990 11836 639882
rect 11796 580984 11848 580990
rect 11796 580926 11848 580932
rect 14476 516118 14504 641038
rect 15844 640892 15896 640898
rect 15844 640834 15896 640840
rect 14556 639872 14608 639878
rect 14556 639814 14608 639820
rect 14568 528562 14596 639814
rect 14556 528556 14608 528562
rect 14556 528498 14608 528504
rect 14464 516112 14516 516118
rect 14464 516054 14516 516060
rect 15856 463690 15884 640834
rect 18604 640416 18656 640422
rect 18604 640358 18656 640364
rect 15936 639804 15988 639810
rect 15936 639746 15988 639752
rect 15948 476066 15976 639746
rect 17316 639668 17368 639674
rect 17316 639610 17368 639616
rect 17224 638308 17276 638314
rect 17224 638250 17276 638256
rect 15936 476060 15988 476066
rect 15936 476002 15988 476008
rect 15844 463684 15896 463690
rect 15844 463626 15896 463632
rect 17236 411262 17264 638250
rect 17328 423638 17356 639610
rect 17316 423632 17368 423638
rect 17316 423574 17368 423580
rect 17224 411256 17276 411262
rect 17224 411198 17276 411204
rect 18616 255270 18644 640358
rect 18696 639600 18748 639606
rect 18696 639542 18748 639548
rect 18708 372570 18736 639542
rect 21456 639464 21508 639470
rect 21456 639406 21508 639412
rect 21364 637628 21416 637634
rect 21364 637570 21416 637576
rect 18696 372564 18748 372570
rect 18696 372506 18748 372512
rect 18604 255264 18656 255270
rect 18604 255206 18656 255212
rect 21376 97986 21404 637570
rect 21468 320142 21496 639406
rect 22744 639396 22796 639402
rect 22744 639338 22796 639344
rect 21456 320136 21508 320142
rect 21456 320078 21508 320084
rect 22756 267714 22784 639338
rect 25504 639260 25556 639266
rect 25504 639202 25556 639208
rect 22744 267708 22796 267714
rect 22744 267650 22796 267656
rect 25516 215286 25544 639202
rect 29642 639160 29698 639169
rect 29642 639095 29698 639104
rect 25504 215280 25556 215286
rect 25504 215222 25556 215228
rect 21364 97980 21416 97986
rect 21364 97922 21416 97928
rect 11704 85536 11756 85542
rect 11704 85478 11756 85484
rect 23388 63504 23440 63510
rect 23388 63446 23440 63452
rect 20628 63300 20680 63306
rect 20628 63242 20680 63248
rect 10968 63232 11020 63238
rect 10968 63174 11020 63180
rect 6828 62892 6880 62898
rect 6828 62834 6880 62840
rect 4896 61464 4948 61470
rect 4896 61406 4948 61412
rect 4804 58948 4856 58954
rect 4804 58890 4856 58896
rect 4908 3534 4936 61406
rect 6840 6914 6868 62834
rect 8208 61396 8260 61402
rect 8208 61338 8260 61344
rect 6472 6886 6868 6914
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6472 480 6500 6886
rect 8220 3534 8248 61338
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7668 480 7696 3470
rect 8772 480 8800 3538
rect 10980 3534 11008 63174
rect 12348 63164 12400 63170
rect 12348 63106 12400 63112
rect 12256 3868 12308 3874
rect 12256 3810 12308 3816
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12268 1986 12296 3810
rect 12360 3534 12388 63106
rect 16488 63028 16540 63034
rect 16488 62970 16540 62976
rect 13728 62960 13780 62966
rect 13728 62902 13780 62908
rect 13740 6914 13768 62902
rect 15108 62280 15160 62286
rect 15108 62222 15160 62228
rect 15120 6914 15148 62222
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12268 1958 12388 1986
rect 12360 480 12388 1958
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3602 16528 62970
rect 18604 61736 18656 61742
rect 18604 61678 18656 61684
rect 17868 61532 17920 61538
rect 17868 61474 17920 61480
rect 17880 3602 17908 61474
rect 18616 3670 18644 61678
rect 20536 3800 20588 3806
rect 20536 3742 20588 3748
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 15948 480 15976 3538
rect 17052 480 17080 3538
rect 18248 480 18276 3538
rect 19444 480 19472 3538
rect 20548 1986 20576 3742
rect 20640 3602 20668 63242
rect 22008 61600 22060 61606
rect 22008 61542 22060 61548
rect 22020 6914 22048 61542
rect 23400 6914 23428 63446
rect 24768 63436 24820 63442
rect 24768 63378 24820 63384
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20548 1958 20668 1986
rect 20640 480 20668 1958
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3602 24808 63378
rect 26148 63368 26200 63374
rect 26148 63310 26200 63316
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24228 480 24256 3538
rect 26160 3398 26188 63310
rect 29656 33114 29684 639095
rect 32416 137970 32444 641650
rect 176936 641640 176988 641646
rect 176936 641582 176988 641588
rect 43536 641572 43588 641578
rect 43536 641514 43588 641520
rect 40684 640960 40736 640966
rect 40684 640902 40736 640908
rect 33782 640656 33838 640665
rect 33782 640591 33838 640600
rect 32494 636304 32550 636313
rect 32494 636239 32550 636248
rect 32508 607170 32536 636239
rect 32496 607164 32548 607170
rect 32496 607106 32548 607112
rect 32404 137964 32456 137970
rect 32404 137906 32456 137912
rect 33048 62756 33100 62762
rect 33048 62698 33100 62704
rect 29736 61940 29788 61946
rect 29736 61882 29788 61888
rect 29644 33108 29696 33114
rect 29644 33050 29696 33056
rect 29748 3874 29776 61882
rect 30104 4820 30156 4826
rect 30104 4762 30156 4768
rect 29736 3868 29788 3874
rect 29736 3810 29788 3816
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 25332 480 25360 3334
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26528 480 26556 3130
rect 27724 480 27752 3334
rect 28908 3324 28960 3330
rect 28908 3266 28960 3272
rect 28920 480 28948 3266
rect 30116 480 30144 4762
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31312 480 31340 4014
rect 33060 3602 33088 62698
rect 33796 45558 33824 640591
rect 36544 639192 36596 639198
rect 36544 639134 36596 639140
rect 35164 636880 35216 636886
rect 35164 636822 35216 636828
rect 33874 636440 33930 636449
rect 33874 636375 33930 636384
rect 33888 554742 33916 636375
rect 33876 554736 33928 554742
rect 33876 554678 33928 554684
rect 34428 62620 34480 62626
rect 34428 62562 34480 62568
rect 33784 45552 33836 45558
rect 33784 45494 33836 45500
rect 34440 3602 34468 62562
rect 35176 6866 35204 636822
rect 35254 636712 35310 636721
rect 35254 636647 35310 636656
rect 35268 502314 35296 636647
rect 35256 502308 35308 502314
rect 35256 502250 35308 502256
rect 36556 164218 36584 639134
rect 39304 639124 39356 639130
rect 39304 639066 39356 639072
rect 36544 164212 36596 164218
rect 36544 164154 36596 164160
rect 39316 111790 39344 639066
rect 40696 358766 40724 640902
rect 40868 638784 40920 638790
rect 40868 638726 40920 638732
rect 40774 637392 40830 637401
rect 40774 637327 40830 637336
rect 40788 449886 40816 637327
rect 40880 619614 40908 638726
rect 43444 638444 43496 638450
rect 43444 638386 43496 638392
rect 40868 619608 40920 619614
rect 40868 619550 40920 619556
rect 40776 449880 40828 449886
rect 40776 449822 40828 449828
rect 40684 358760 40736 358766
rect 40684 358702 40736 358708
rect 43456 293962 43484 638386
rect 43548 567186 43576 641514
rect 139400 641368 139452 641374
rect 139400 641310 139452 641316
rect 50436 641300 50488 641306
rect 50436 641242 50488 641248
rect 50344 640824 50396 640830
rect 50344 640766 50396 640772
rect 47584 639056 47636 639062
rect 47584 638998 47636 639004
rect 43536 567180 43588 567186
rect 43536 567122 43588 567128
rect 43444 293956 43496 293962
rect 43444 293898 43496 293904
rect 39304 111784 39356 111790
rect 39304 111726 39356 111732
rect 47596 71738 47624 638998
rect 50356 306338 50384 640766
rect 50448 398818 50476 641242
rect 53196 641232 53248 641238
rect 53196 641174 53248 641180
rect 51724 640688 51776 640694
rect 51724 640630 51776 640636
rect 50436 398812 50488 398818
rect 50436 398754 50488 398760
rect 50344 306332 50396 306338
rect 50344 306274 50396 306280
rect 51736 241466 51764 640630
rect 53104 640484 53156 640490
rect 53104 640426 53156 640432
rect 51724 241460 51776 241466
rect 51724 241402 51776 241408
rect 53116 150414 53144 640426
rect 53208 346390 53236 641174
rect 118516 640620 118568 640626
rect 118516 640562 118568 640568
rect 105912 640552 105964 640558
rect 72514 640520 72570 640529
rect 105912 640494 105964 640500
rect 72514 640455 72570 640464
rect 68374 639296 68430 639305
rect 68374 639231 68430 639240
rect 55862 639024 55918 639033
rect 55862 638959 55918 638968
rect 55876 638452 55904 638959
rect 68388 638452 68416 639231
rect 72528 638452 72556 640455
rect 93400 639328 93452 639334
rect 93400 639270 93452 639276
rect 80888 638988 80940 638994
rect 80888 638930 80940 638936
rect 80900 638452 80928 638930
rect 93412 638452 93440 639270
rect 105924 638452 105952 640494
rect 118528 638452 118556 640562
rect 131028 639532 131080 639538
rect 131028 639474 131080 639480
rect 131040 638452 131068 639474
rect 139412 638452 139440 641310
rect 168564 641164 168616 641170
rect 168564 641106 168616 641112
rect 143540 640756 143592 640762
rect 143540 640698 143592 640704
rect 143552 638452 143580 640698
rect 164424 640348 164476 640354
rect 164424 640290 164476 640296
rect 156052 639736 156104 639742
rect 156052 639678 156104 639684
rect 152280 638512 152332 638518
rect 151938 638460 152280 638466
rect 151938 638454 152332 638460
rect 151938 638438 152320 638454
rect 156064 638452 156092 639678
rect 160560 638580 160612 638586
rect 160560 638522 160612 638528
rect 160572 638466 160600 638522
rect 160310 638438 160600 638466
rect 164436 638452 164464 640290
rect 168576 638452 168604 641106
rect 172796 641028 172848 641034
rect 172796 640970 172848 640976
rect 172808 638452 172836 640970
rect 175924 640348 175976 640354
rect 175924 640290 175976 640296
rect 175936 638722 175964 640290
rect 175924 638716 175976 638722
rect 175924 638658 175976 638664
rect 176948 638452 176976 641582
rect 189448 641504 189500 641510
rect 189448 641446 189500 641452
rect 189080 641368 189132 641374
rect 189080 641310 189132 641316
rect 181168 640076 181220 640082
rect 181168 640018 181220 640024
rect 181180 638452 181208 640018
rect 189092 638858 189120 641310
rect 189080 638852 189132 638858
rect 189080 638794 189132 638800
rect 189460 638452 189488 641446
rect 214564 641436 214616 641442
rect 214564 641378 214616 641384
rect 202052 641368 202104 641374
rect 202052 641310 202104 641316
rect 193680 640144 193732 640150
rect 193680 640086 193732 640092
rect 193692 638452 193720 640086
rect 202064 638452 202092 641310
rect 206192 640212 206244 640218
rect 206192 640154 206244 640160
rect 206204 638452 206232 640154
rect 214576 638452 214604 641378
rect 218704 640280 218756 640286
rect 218704 640222 218756 640228
rect 218716 638452 218744 640222
rect 222948 638452 222976 643078
rect 227076 638920 227128 638926
rect 227076 638862 227128 638868
rect 227088 638452 227116 638862
rect 231688 638466 231716 644446
rect 235920 638466 235948 696934
rect 240048 683256 240100 683262
rect 240048 683198 240100 683204
rect 240060 644474 240088 683198
rect 242176 668642 242204 700470
rect 242164 668636 242216 668642
rect 242164 668578 242216 668584
rect 239968 644446 240088 644474
rect 239968 638466 239996 644446
rect 243820 642388 243872 642394
rect 243820 642330 243872 642336
rect 231242 638438 231716 638466
rect 235474 638438 235948 638466
rect 239614 638438 239996 638466
rect 243832 638452 243860 642330
rect 248340 638466 248368 700538
rect 252468 700528 252520 700534
rect 252468 700470 252520 700476
rect 252480 638466 252508 700470
rect 256332 643748 256384 643754
rect 256332 643690 256384 643696
rect 247986 638438 248368 638466
rect 252126 638438 252508 638466
rect 256344 638452 256372 643690
rect 260760 638466 260788 700810
rect 264888 700800 264940 700806
rect 264888 700742 264940 700748
rect 264900 638466 264928 700742
rect 267660 699854 267688 703520
rect 277308 700256 277360 700262
rect 277308 700198 277360 700204
rect 273168 700188 273220 700194
rect 273168 700130 273220 700136
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 268844 642592 268896 642598
rect 268844 642534 268896 642540
rect 260498 638438 260788 638466
rect 264730 638438 264928 638466
rect 268856 638452 268884 642534
rect 273180 638466 273208 700130
rect 277320 638466 277348 700198
rect 283852 699786 283880 703520
rect 289728 699984 289780 699990
rect 289728 699926 289780 699932
rect 285588 699916 285640 699922
rect 285588 699858 285640 699864
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 281356 642660 281408 642666
rect 281356 642602 281408 642608
rect 273010 638438 273208 638466
rect 277242 638438 277348 638466
rect 281368 638452 281396 642602
rect 285600 638452 285628 699858
rect 289740 638452 289768 699926
rect 298100 699848 298152 699854
rect 298100 699790 298152 699796
rect 293960 642728 294012 642734
rect 293960 642670 294012 642676
rect 293972 638452 294000 642670
rect 298112 638452 298140 699790
rect 299492 642734 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 327080 701004 327132 701010
rect 327080 700946 327132 700952
rect 322940 700936 322992 700942
rect 322940 700878 322992 700884
rect 310520 700120 310572 700126
rect 310520 700062 310572 700068
rect 302240 699780 302292 699786
rect 302240 699722 302292 699728
rect 299480 642728 299532 642734
rect 299480 642670 299532 642676
rect 302252 638452 302280 699722
rect 306380 668636 306432 668642
rect 306380 668578 306432 668584
rect 306392 638466 306420 668578
rect 310532 638466 310560 700062
rect 314660 700052 314712 700058
rect 314660 699994 314712 700000
rect 314672 638466 314700 699994
rect 318984 642524 319036 642530
rect 318984 642466 319036 642472
rect 306392 638438 306498 638466
rect 310532 638438 310638 638466
rect 314672 638438 314870 638466
rect 318996 638452 319024 642466
rect 322952 638466 322980 700878
rect 327092 638466 327120 700946
rect 332520 699922 332548 703520
rect 339500 700732 339552 700738
rect 339500 700674 339552 700680
rect 335360 700664 335412 700670
rect 335360 700606 335412 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 331496 642456 331548 642462
rect 331496 642398 331548 642404
rect 322952 638438 323150 638466
rect 327092 638438 327382 638466
rect 331508 638452 331536 642398
rect 335372 638466 335400 700606
rect 339512 638466 339540 700674
rect 342904 700664 342956 700670
rect 342904 700606 342956 700612
rect 342916 642666 342944 700606
rect 343640 700460 343692 700466
rect 343640 700402 343692 700408
rect 342904 642660 342956 642666
rect 342904 642602 342956 642608
rect 343652 638466 343680 700402
rect 347872 700324 347924 700330
rect 347872 700266 347924 700272
rect 347884 638466 347912 700266
rect 348804 699990 348832 703520
rect 364996 700670 365024 703520
rect 364984 700664 365036 700670
rect 364984 700606 365036 700612
rect 351920 700392 351972 700398
rect 351920 700334 351972 700340
rect 349804 700324 349856 700330
rect 349804 700266 349856 700272
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 349816 642598 349844 700266
rect 349804 642592 349856 642598
rect 349804 642534 349856 642540
rect 351932 638466 351960 700334
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 700330 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700330 494836 703520
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 559668 700330 559696 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 457444 700324 457496 700330
rect 457444 700266 457496 700272
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 526444 700324 526496 700330
rect 526444 700266 526496 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 356060 683188 356112 683194
rect 356060 683130 356112 683136
rect 356072 654134 356100 683130
rect 364340 670744 364392 670750
rect 364340 670686 364392 670692
rect 360200 656940 360252 656946
rect 360200 656882 360252 656888
rect 360212 654134 360240 656882
rect 364352 654134 364380 670686
rect 356072 654106 356192 654134
rect 360212 654106 360424 654134
rect 364352 654106 364472 654134
rect 356164 638466 356192 654106
rect 360396 638466 360424 654106
rect 364444 638466 364472 654106
rect 457456 643754 457484 700266
rect 457444 643748 457496 643754
rect 457444 643690 457496 643696
rect 526456 642394 526484 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 526444 642388 526496 642394
rect 526444 642330 526496 642336
rect 486056 641708 486108 641714
rect 486056 641650 486108 641656
rect 369860 641640 369912 641646
rect 369860 641582 369912 641588
rect 369872 640014 369900 641582
rect 390008 641572 390060 641578
rect 390008 641514 390060 641520
rect 369124 640008 369176 640014
rect 369124 639950 369176 639956
rect 369860 640008 369912 640014
rect 369860 639950 369912 639956
rect 335372 638438 335754 638466
rect 339512 638438 339894 638466
rect 343652 638438 344034 638466
rect 347884 638438 348266 638466
rect 351932 638438 352406 638466
rect 356164 638438 356638 638466
rect 360396 638438 360778 638466
rect 364444 638438 364918 638466
rect 369136 638452 369164 639950
rect 381636 639940 381688 639946
rect 381636 639882 381688 639888
rect 377496 638784 377548 638790
rect 377496 638726 377548 638732
rect 377508 638452 377536 638726
rect 381648 638452 381676 639882
rect 390020 638452 390048 641514
rect 423404 641300 423456 641306
rect 423404 641242 423456 641248
rect 402520 641096 402572 641102
rect 402520 641038 402572 641044
rect 415860 641096 415912 641102
rect 415860 641038 415912 641044
rect 394148 639872 394200 639878
rect 394148 639814 394200 639820
rect 394160 638452 394188 639814
rect 402532 638452 402560 641038
rect 415032 640892 415084 640898
rect 415032 640834 415084 640840
rect 406660 639804 406712 639810
rect 406660 639746 406712 639752
rect 406672 638452 406700 639746
rect 415044 638452 415072 640834
rect 415872 638654 415900 641038
rect 419264 639668 419316 639674
rect 419264 639610 419316 639616
rect 415860 638648 415912 638654
rect 415860 638590 415912 638596
rect 419276 638452 419304 639610
rect 423416 638452 423444 641242
rect 435916 641232 435968 641238
rect 435916 641174 435968 641180
rect 435364 640892 435416 640898
rect 435364 640834 435416 640840
rect 431776 639600 431828 639606
rect 431776 639542 431828 639548
rect 431788 638452 431816 639542
rect 135260 638376 135312 638382
rect 135194 638324 135260 638330
rect 135194 638318 135312 638324
rect 135194 638302 135300 638318
rect 427280 638314 427570 638330
rect 427268 638308 427570 638314
rect 427320 638302 427570 638308
rect 427268 638250 427320 638256
rect 148048 638240 148100 638246
rect 126822 638178 126928 638194
rect 147706 638188 148048 638194
rect 435376 638217 435404 640834
rect 435928 638452 435956 641174
rect 477684 641096 477736 641102
rect 477684 641038 477736 641044
rect 440148 640960 440200 640966
rect 440148 640902 440200 640908
rect 440160 638452 440188 640902
rect 452660 640824 452712 640830
rect 452660 640766 452712 640772
rect 444288 639464 444340 639470
rect 444288 639406 444340 639412
rect 444300 638452 444328 639406
rect 448072 638450 448454 638466
rect 452672 638452 452700 640766
rect 461032 640688 461084 640694
rect 461032 640630 461084 640636
rect 456800 639396 456852 639402
rect 456800 639338 456852 639344
rect 456812 638452 456840 639338
rect 461044 638452 461072 640630
rect 465172 640416 465224 640422
rect 465172 640358 465224 640364
rect 465184 638452 465212 640358
rect 469312 639260 469364 639266
rect 469312 639202 469364 639208
rect 469324 638452 469352 639202
rect 477696 638452 477724 641038
rect 481916 639192 481968 639198
rect 481916 639134 481968 639140
rect 481928 638452 481956 639134
rect 486068 638452 486096 641650
rect 536104 641504 536156 641510
rect 536104 641446 536156 641452
rect 527824 640892 527876 640898
rect 527824 640834 527876 640840
rect 515310 640792 515366 640801
rect 515310 640727 515366 640736
rect 511078 640656 511134 640665
rect 511078 640591 511134 640600
rect 490196 640484 490248 640490
rect 490196 640426 490248 640432
rect 490208 638452 490236 640426
rect 494428 639124 494480 639130
rect 494428 639066 494480 639072
rect 494440 638452 494468 639066
rect 506940 639056 506992 639062
rect 506940 638998 506992 639004
rect 506952 638452 506980 638998
rect 511092 638452 511120 640591
rect 515324 638452 515352 640727
rect 519450 639160 519506 639169
rect 519450 639095 519506 639104
rect 519464 638452 519492 639095
rect 527836 638452 527864 640834
rect 531964 640552 532016 640558
rect 531964 640494 532016 640500
rect 530584 639328 530636 639334
rect 530584 639270 530636 639276
rect 448060 638444 448454 638450
rect 448112 638438 448454 638444
rect 448060 638386 448112 638392
rect 473372 638314 473570 638330
rect 502536 638314 502826 638330
rect 523328 638314 523710 638330
rect 473360 638308 473570 638314
rect 473412 638302 473570 638308
rect 502524 638308 502826 638314
rect 473360 638250 473412 638256
rect 502576 638302 502826 638308
rect 523316 638308 523710 638314
rect 502524 638250 502576 638256
rect 523368 638302 523710 638308
rect 523316 638250 523368 638256
rect 147706 638182 148100 638188
rect 435362 638208 435418 638217
rect 126822 638172 126940 638178
rect 126822 638166 126888 638172
rect 147706 638166 148088 638182
rect 435362 638143 435418 638152
rect 126888 638114 126940 638120
rect 114468 638104 114520 638110
rect 101798 638042 102088 638058
rect 114310 638052 114468 638058
rect 114310 638046 114520 638052
rect 101798 638036 102100 638042
rect 101798 638030 102048 638036
rect 114310 638030 114508 638046
rect 102048 637978 102100 637984
rect 97908 637968 97960 637974
rect 60186 637936 60242 637945
rect 60030 637894 60186 637922
rect 64418 637936 64474 637945
rect 64170 637894 64418 637922
rect 60186 637871 60242 637880
rect 77022 637936 77078 637945
rect 76774 637894 77022 637922
rect 64418 637871 64474 637880
rect 85210 637936 85266 637945
rect 85054 637894 85210 637922
rect 77022 637871 77078 637880
rect 89286 637906 89576 637922
rect 97658 637916 97908 637922
rect 110328 637968 110380 637974
rect 97658 637910 97960 637916
rect 110170 637916 110328 637922
rect 122748 637968 122800 637974
rect 110170 637910 110380 637916
rect 122682 637916 122748 637922
rect 185490 637936 185546 637945
rect 122682 637910 122800 637916
rect 89286 637900 89588 637906
rect 89286 637894 89536 637900
rect 85210 637871 85266 637880
rect 97658 637894 97948 637910
rect 110170 637894 110368 637910
rect 122682 637894 122788 637910
rect 185334 637894 185490 637922
rect 198002 637936 198058 637945
rect 197846 637894 198002 637922
rect 185490 637871 185546 637880
rect 210514 637936 210570 637945
rect 210358 637894 210514 637922
rect 198002 637871 198058 637880
rect 210514 637871 210570 637880
rect 373078 637936 373134 637945
rect 385590 637936 385646 637945
rect 373134 637894 373290 637922
rect 373078 637871 373134 637880
rect 398102 637936 398158 637945
rect 385646 637894 385802 637922
rect 385590 637871 385646 637880
rect 410614 637936 410670 637945
rect 398158 637894 398406 637922
rect 398102 637871 398158 637880
rect 498290 637936 498346 637945
rect 410670 637894 410918 637922
rect 410614 637871 410670 637880
rect 498346 637894 498594 637922
rect 498290 637871 498346 637880
rect 89536 637842 89588 637848
rect 53196 346384 53248 346390
rect 53196 346326 53248 346332
rect 53104 150408 53156 150414
rect 53104 150350 53156 150356
rect 530596 126954 530624 639270
rect 530676 638920 530728 638926
rect 530676 638862 530728 638868
rect 530688 632058 530716 638862
rect 530676 632052 530728 632058
rect 530676 631994 530728 632000
rect 531976 167006 532004 640494
rect 533436 640076 533488 640082
rect 533436 640018 533488 640024
rect 532056 638512 532108 638518
rect 532056 638454 532108 638460
rect 532068 313274 532096 638454
rect 533342 637800 533398 637809
rect 533342 637735 533398 637744
rect 532056 313268 532108 313274
rect 532056 313210 532108 313216
rect 531964 167000 532016 167006
rect 531964 166942 532016 166948
rect 530584 126948 530636 126954
rect 530584 126890 530636 126896
rect 47584 71732 47636 71738
rect 47584 71674 47636 71680
rect 39948 62688 40000 62694
rect 39948 62630 40000 62636
rect 36544 62008 36596 62014
rect 36544 61950 36596 61956
rect 35256 61872 35308 61878
rect 35256 61814 35308 61820
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 34796 3868 34848 3874
rect 34796 3810 34848 3816
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 32416 480 32444 3538
rect 33612 480 33640 3538
rect 34808 480 34836 3810
rect 35268 3194 35296 61814
rect 36556 3738 36584 61950
rect 39960 6914 39988 62630
rect 41328 62552 41380 62558
rect 41328 62494 41380 62500
rect 39592 6886 39988 6914
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 35992 3256 36044 3262
rect 35992 3198 36044 3204
rect 35256 3188 35308 3194
rect 35256 3130 35308 3136
rect 36004 480 36032 3198
rect 37188 3188 37240 3194
rect 37188 3130 37240 3136
rect 37200 480 37228 3130
rect 38396 480 38424 3878
rect 39592 480 39620 6886
rect 41340 3398 41368 62494
rect 50988 62484 51040 62490
rect 50988 62426 51040 62432
rect 43444 62416 43496 62422
rect 43444 62358 43496 62364
rect 43456 4078 43484 62358
rect 48228 61668 48280 61674
rect 48228 61610 48280 61616
rect 48240 6914 48268 61610
rect 47872 6886 48268 6914
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 43444 4072 43496 4078
rect 43444 4014 43496 4020
rect 41880 4004 41932 4010
rect 41880 3946 41932 3952
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3946
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 43088 480 43116 3334
rect 44272 3052 44324 3058
rect 44272 2994 44324 3000
rect 44284 480 44312 2994
rect 45480 480 45508 4082
rect 46664 2984 46716 2990
rect 46664 2926 46716 2932
rect 46676 480 46704 2926
rect 47872 480 47900 6886
rect 51000 3738 51028 62426
rect 53104 62348 53156 62354
rect 53104 62290 53156 62296
rect 52368 61804 52420 61810
rect 52368 61746 52420 61752
rect 52380 3738 52408 61746
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 50988 3732 51040 3738
rect 50988 3674 51040 3680
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 52368 3732 52420 3738
rect 52368 3674 52420 3680
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48976 480 49004 3130
rect 50172 480 50200 3674
rect 51368 480 51396 3674
rect 53116 3194 53144 62290
rect 54312 61742 54340 65484
rect 55232 62014 55260 65484
rect 55864 62212 55916 62218
rect 55864 62154 55916 62160
rect 55220 62008 55272 62014
rect 55220 61950 55272 61956
rect 54300 61736 54352 61742
rect 54300 61678 54352 61684
rect 55128 61736 55180 61742
rect 55128 61678 55180 61684
rect 55140 6914 55168 61678
rect 54956 6886 55168 6914
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 53104 3188 53156 3194
rect 53104 3130 53156 3136
rect 52552 2916 52604 2922
rect 52552 2858 52604 2864
rect 52564 480 52592 2858
rect 53760 480 53788 4014
rect 54956 480 54984 6886
rect 55876 3126 55904 62154
rect 56152 61470 56180 65484
rect 57164 62830 57192 65484
rect 57152 62824 57204 62830
rect 57152 62766 57204 62772
rect 57888 62824 57940 62830
rect 57888 62766 57940 62772
rect 56140 61464 56192 61470
rect 56140 61406 56192 61412
rect 57900 3534 57928 62766
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 55864 3120 55916 3126
rect 55864 3062 55916 3068
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 56060 480 56088 2926
rect 57256 480 57284 3470
rect 58084 3466 58112 65484
rect 59096 62898 59124 65484
rect 60016 64874 60044 65484
rect 59924 64846 60044 64874
rect 59084 62892 59136 62898
rect 59084 62834 59136 62840
rect 59924 61402 59952 64846
rect 61028 62150 61056 65484
rect 61948 63238 61976 65484
rect 61936 63232 61988 63238
rect 61936 63174 61988 63180
rect 62960 63170 62988 65484
rect 62948 63164 63000 63170
rect 62948 63106 63000 63112
rect 62764 62892 62816 62898
rect 62764 62834 62816 62840
rect 60004 62144 60056 62150
rect 60004 62086 60056 62092
rect 61016 62144 61068 62150
rect 61016 62086 61068 62092
rect 61384 62144 61436 62150
rect 61384 62086 61436 62092
rect 59912 61396 59964 61402
rect 59912 61338 59964 61344
rect 58440 6180 58492 6186
rect 58440 6122 58492 6128
rect 58072 3460 58124 3466
rect 58072 3402 58124 3408
rect 58452 480 58480 6122
rect 60016 3330 60044 62086
rect 60832 3460 60884 3466
rect 60832 3402 60884 3408
rect 60004 3324 60056 3330
rect 60004 3266 60056 3272
rect 59636 2848 59688 2854
rect 59636 2790 59688 2796
rect 59648 480 59676 2790
rect 60844 480 60872 3402
rect 61396 3262 61424 62086
rect 62028 4888 62080 4894
rect 62028 4830 62080 4836
rect 61384 3256 61436 3262
rect 61384 3198 61436 3204
rect 62040 480 62068 4830
rect 62776 3806 62804 62834
rect 63880 61946 63908 65484
rect 64144 63164 64196 63170
rect 64144 63106 64196 63112
rect 63868 61940 63920 61946
rect 63868 61882 63920 61888
rect 62764 3800 62816 3806
rect 62764 3742 62816 3748
rect 64156 3262 64184 63106
rect 64892 62966 64920 65484
rect 65524 63096 65576 63102
rect 65524 63038 65576 63044
rect 64880 62960 64932 62966
rect 64880 62902 64932 62908
rect 65536 6914 65564 63038
rect 65812 62286 65840 65484
rect 66824 63034 66852 65484
rect 66812 63028 66864 63034
rect 66812 62970 66864 62976
rect 65800 62280 65852 62286
rect 65800 62222 65852 62228
rect 66904 62280 66956 62286
rect 66904 62222 66956 62228
rect 66168 61396 66220 61402
rect 66168 61338 66220 61344
rect 65444 6886 65564 6914
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64144 3256 64196 3262
rect 64144 3198 64196 3204
rect 63224 3120 63276 3126
rect 63224 3062 63276 3068
rect 63236 480 63264 3062
rect 64340 480 64368 3470
rect 65444 3058 65472 6886
rect 66180 3602 66208 61338
rect 65524 3596 65576 3602
rect 65524 3538 65576 3544
rect 66168 3596 66220 3602
rect 66168 3538 66220 3544
rect 65432 3052 65484 3058
rect 65432 2994 65484 3000
rect 65536 480 65564 3538
rect 66720 3256 66772 3262
rect 66720 3198 66772 3204
rect 66732 480 66760 3198
rect 66916 2922 66944 62222
rect 67744 61538 67772 65484
rect 67732 61532 67784 61538
rect 67732 61474 67784 61480
rect 68756 3670 68784 65484
rect 69676 63306 69704 65484
rect 69664 63300 69716 63306
rect 69664 63242 69716 63248
rect 70688 62898 70716 65484
rect 70676 62892 70728 62898
rect 70676 62834 70728 62840
rect 71608 61606 71636 65484
rect 72620 63510 72648 65484
rect 72608 63504 72660 63510
rect 72608 63446 72660 63452
rect 73540 63442 73568 65484
rect 73528 63436 73580 63442
rect 73528 63378 73580 63384
rect 74552 63374 74580 65484
rect 74540 63368 74592 63374
rect 74540 63310 74592 63316
rect 75276 63368 75328 63374
rect 75276 63310 75328 63316
rect 72424 63028 72476 63034
rect 72424 62970 72476 62976
rect 71688 62960 71740 62966
rect 71688 62902 71740 62908
rect 71596 61600 71648 61606
rect 71596 61542 71648 61548
rect 70308 61532 70360 61538
rect 70308 61474 70360 61480
rect 68744 3664 68796 3670
rect 68744 3606 68796 3612
rect 70320 3602 70348 61474
rect 71700 6914 71728 62902
rect 71516 6886 71728 6914
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 67916 3052 67968 3058
rect 67916 2994 67968 3000
rect 66904 2916 66956 2922
rect 66904 2858 66956 2864
rect 67928 480 67956 2994
rect 69124 480 69152 3538
rect 70308 3324 70360 3330
rect 70308 3266 70360 3272
rect 70320 480 70348 3266
rect 71516 480 71544 6886
rect 72436 4826 72464 62970
rect 73804 62892 73856 62898
rect 73804 62834 73856 62840
rect 73068 61464 73120 61470
rect 73068 61406 73120 61412
rect 72424 4820 72476 4826
rect 72424 4762 72476 4768
rect 73080 3602 73108 61406
rect 73816 3670 73844 62834
rect 75184 62144 75236 62150
rect 75184 62086 75236 62092
rect 75196 3874 75224 62086
rect 75184 3868 75236 3874
rect 75184 3810 75236 3816
rect 73804 3664 73856 3670
rect 73804 3606 73856 3612
rect 75000 3664 75052 3670
rect 75000 3606 75052 3612
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 72620 480 72648 3538
rect 73804 3052 73856 3058
rect 73804 2994 73856 3000
rect 73816 480 73844 2994
rect 75012 480 75040 3606
rect 75288 2922 75316 63310
rect 75472 61878 75500 65484
rect 76484 62898 76512 65484
rect 77404 63238 77432 65484
rect 77392 63232 77444 63238
rect 77392 63174 77444 63180
rect 77944 63232 77996 63238
rect 77944 63174 77996 63180
rect 76472 62892 76524 62898
rect 76472 62834 76524 62840
rect 76564 62892 76616 62898
rect 76564 62834 76616 62840
rect 75460 61872 75512 61878
rect 75460 61814 75512 61820
rect 76576 3806 76604 62834
rect 77208 61600 77260 61606
rect 77208 61542 77260 61548
rect 76564 3800 76616 3806
rect 76564 3742 76616 3748
rect 77220 3602 77248 61542
rect 77392 3936 77444 3942
rect 77392 3878 77444 3884
rect 76196 3596 76248 3602
rect 76196 3538 76248 3544
rect 77208 3596 77260 3602
rect 77208 3538 77260 3544
rect 75276 2916 75328 2922
rect 75276 2858 75328 2864
rect 76208 480 76236 3538
rect 77404 480 77432 3878
rect 77956 3398 77984 63174
rect 78416 63034 78444 65484
rect 78404 63028 78456 63034
rect 78404 62970 78456 62976
rect 79336 62422 79364 65484
rect 79416 63300 79468 63306
rect 79416 63242 79468 63248
rect 79324 62416 79376 62422
rect 79324 62358 79376 62364
rect 79428 45554 79456 63242
rect 80348 62762 80376 65484
rect 80336 62756 80388 62762
rect 80336 62698 80388 62704
rect 80704 62756 80756 62762
rect 80704 62698 80756 62704
rect 79968 61872 80020 61878
rect 79968 61814 80020 61820
rect 79336 45526 79456 45554
rect 79336 4010 79364 45526
rect 79980 6914 80008 61814
rect 79704 6886 80008 6914
rect 79324 4004 79376 4010
rect 79324 3946 79376 3952
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 77944 3392 77996 3398
rect 77944 3334 77996 3340
rect 78600 480 78628 3810
rect 79704 480 79732 6886
rect 80716 4146 80744 62698
rect 81268 62626 81296 65484
rect 81348 63028 81400 63034
rect 81348 62970 81400 62976
rect 81256 62620 81308 62626
rect 81256 62562 81308 62568
rect 80704 4140 80756 4146
rect 80704 4082 80756 4088
rect 81360 3602 81388 62970
rect 82280 62150 82308 65484
rect 83200 63170 83228 65484
rect 83188 63164 83240 63170
rect 83188 63106 83240 63112
rect 84212 62218 84240 65484
rect 84844 63504 84896 63510
rect 84844 63446 84896 63452
rect 84200 62212 84252 62218
rect 84200 62154 84252 62160
rect 82268 62144 82320 62150
rect 82268 62086 82320 62092
rect 84108 61940 84160 61946
rect 84108 61882 84160 61888
rect 80888 3596 80940 3602
rect 80888 3538 80940 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 82084 3596 82136 3602
rect 82084 3538 82136 3544
rect 80900 480 80928 3538
rect 82096 480 82124 3538
rect 84120 3398 84148 61882
rect 83280 3392 83332 3398
rect 83280 3334 83332 3340
rect 84108 3392 84160 3398
rect 84108 3334 84160 3340
rect 83292 480 83320 3334
rect 84856 3194 84884 63446
rect 85132 62966 85160 65484
rect 85120 62960 85172 62966
rect 85120 62902 85172 62908
rect 86144 62694 86172 65484
rect 86868 63164 86920 63170
rect 86868 63106 86920 63112
rect 86132 62688 86184 62694
rect 86132 62630 86184 62636
rect 86776 6248 86828 6254
rect 86776 6190 86828 6196
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 84844 3188 84896 3194
rect 84844 3130 84896 3136
rect 84476 2916 84528 2922
rect 84476 2858 84528 2864
rect 84488 480 84516 2858
rect 85684 480 85712 3334
rect 86788 3210 86816 6190
rect 86880 3398 86908 63106
rect 87064 62558 87092 65484
rect 87604 63436 87656 63442
rect 87604 63378 87656 63384
rect 87052 62552 87104 62558
rect 87052 62494 87104 62500
rect 86868 3392 86920 3398
rect 86868 3334 86920 3340
rect 86788 3182 86908 3210
rect 86880 480 86908 3182
rect 87616 3126 87644 63378
rect 88076 63306 88104 65484
rect 88064 63300 88116 63306
rect 88064 63242 88116 63248
rect 88996 63238 89024 65484
rect 88984 63232 89036 63238
rect 88984 63174 89036 63180
rect 90008 63102 90036 65484
rect 90364 63300 90416 63306
rect 90364 63242 90416 63248
rect 89996 63096 90048 63102
rect 89996 63038 90048 63044
rect 88248 62960 88300 62966
rect 88248 62902 88300 62908
rect 88260 6914 88288 62902
rect 88984 62144 89036 62150
rect 88984 62086 89036 62092
rect 87984 6886 88288 6914
rect 87604 3120 87656 3126
rect 87604 3062 87656 3068
rect 87984 480 88012 6886
rect 88996 3738 89024 62086
rect 90376 6914 90404 63242
rect 90928 62762 90956 65484
rect 90916 62756 90968 62762
rect 90916 62698 90968 62704
rect 91744 62756 91796 62762
rect 91744 62698 91796 62704
rect 91008 62008 91060 62014
rect 91008 61950 91060 61956
rect 90284 6886 90404 6914
rect 90284 4078 90312 6886
rect 90272 4072 90324 4078
rect 90272 4014 90324 4020
rect 89168 4004 89220 4010
rect 89168 3946 89220 3952
rect 88984 3732 89036 3738
rect 88984 3674 89036 3680
rect 89180 480 89208 3946
rect 91020 3398 91048 61950
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 90376 480 90404 3334
rect 91560 3188 91612 3194
rect 91560 3130 91612 3136
rect 91572 480 91600 3130
rect 91756 2990 91784 62698
rect 91940 62150 91968 65484
rect 91928 62144 91980 62150
rect 91928 62086 91980 62092
rect 92860 61674 92888 65484
rect 93768 63232 93820 63238
rect 93768 63174 93820 63180
rect 92848 61668 92900 61674
rect 92848 61610 92900 61616
rect 93780 3262 93808 63174
rect 93872 62354 93900 65484
rect 94792 62490 94820 65484
rect 95148 63096 95200 63102
rect 95148 63038 95200 63044
rect 94780 62484 94832 62490
rect 94780 62426 94832 62432
rect 93860 62348 93912 62354
rect 93860 62290 93912 62296
rect 95056 61668 95108 61674
rect 95056 61610 95108 61616
rect 92756 3256 92808 3262
rect 92756 3198 92808 3204
rect 93768 3256 93820 3262
rect 93768 3198 93820 3204
rect 91744 2984 91796 2990
rect 91744 2926 91796 2932
rect 92768 480 92796 3198
rect 95068 2922 95096 61610
rect 93952 2916 94004 2922
rect 93952 2858 94004 2864
rect 95056 2916 95108 2922
rect 95056 2858 95108 2864
rect 93964 480 93992 2858
rect 95160 480 95188 63038
rect 95804 61810 95832 65484
rect 95884 62552 95936 62558
rect 95884 62494 95936 62500
rect 95792 61804 95844 61810
rect 95792 61746 95844 61752
rect 95896 3330 95924 62494
rect 96724 62286 96752 65484
rect 97736 63306 97764 65484
rect 98656 64874 98684 65484
rect 98564 64846 98684 64874
rect 97724 63300 97776 63306
rect 97724 63242 97776 63248
rect 97264 62620 97316 62626
rect 97264 62562 97316 62568
rect 96712 62280 96764 62286
rect 96712 62222 96764 62228
rect 96252 4072 96304 4078
rect 96252 4014 96304 4020
rect 95884 3324 95936 3330
rect 95884 3266 95936 3272
rect 96264 480 96292 4014
rect 97276 3466 97304 62562
rect 97908 61804 97960 61810
rect 97908 61746 97960 61752
rect 97920 3534 97948 61746
rect 98564 61742 98592 64846
rect 99668 63374 99696 65484
rect 99656 63368 99708 63374
rect 99656 63310 99708 63316
rect 99288 63300 99340 63306
rect 99288 63242 99340 63248
rect 98644 62280 98696 62286
rect 98644 62222 98696 62228
rect 98552 61736 98604 61742
rect 98552 61678 98604 61684
rect 98656 6914 98684 62222
rect 98564 6886 98684 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 97264 3460 97316 3466
rect 97264 3402 97316 3408
rect 97460 480 97488 3470
rect 98564 3058 98592 6886
rect 99300 3534 99328 63242
rect 100588 62830 100616 65484
rect 100576 62824 100628 62830
rect 100576 62766 100628 62772
rect 100116 62484 100168 62490
rect 100116 62426 100168 62432
rect 100024 62144 100076 62150
rect 100024 62086 100076 62092
rect 99840 3936 99892 3942
rect 99840 3878 99892 3884
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 98552 3052 98604 3058
rect 98552 2994 98604 3000
rect 98656 480 98684 3470
rect 99852 480 99880 3878
rect 100036 3262 100064 62086
rect 100128 3738 100156 62426
rect 101600 6186 101628 65484
rect 102520 63510 102548 65484
rect 102508 63504 102560 63510
rect 102508 63446 102560 63452
rect 103428 62824 103480 62830
rect 103428 62766 103480 62772
rect 101588 6180 101640 6186
rect 101588 6122 101640 6128
rect 101036 6112 101088 6118
rect 101036 6054 101088 6060
rect 100116 3732 100168 3738
rect 100116 3674 100168 3680
rect 100024 3256 100076 3262
rect 100024 3198 100076 3204
rect 101048 480 101076 6054
rect 103336 3732 103388 3738
rect 103336 3674 103388 3680
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 102244 480 102272 3470
rect 103348 480 103376 3674
rect 103440 3534 103468 62766
rect 103532 62150 103560 65484
rect 103520 62144 103572 62150
rect 103520 62086 103572 62092
rect 104452 4894 104480 65484
rect 105464 63442 105492 65484
rect 105544 63504 105596 63510
rect 105544 63446 105596 63452
rect 105452 63436 105504 63442
rect 105452 63378 105504 63384
rect 104440 4888 104492 4894
rect 104440 4830 104492 4836
rect 105556 3806 105584 63446
rect 106188 63368 106240 63374
rect 106188 63310 106240 63316
rect 105544 3800 105596 3806
rect 105544 3742 105596 3748
rect 106200 3534 106228 63310
rect 106384 62626 106412 65484
rect 106372 62620 106424 62626
rect 106372 62562 106424 62568
rect 107016 62620 107068 62626
rect 107016 62562 107068 62568
rect 106924 62212 106976 62218
rect 106924 62154 106976 62160
rect 106936 3670 106964 62154
rect 106924 3664 106976 3670
rect 106924 3606 106976 3612
rect 103428 3528 103480 3534
rect 103428 3470 103480 3476
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 104532 3460 104584 3466
rect 104532 3402 104584 3408
rect 104544 480 104572 3402
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 107028 3398 107056 62562
rect 107396 61402 107424 65484
rect 108316 62762 108344 65484
rect 108304 62756 108356 62762
rect 108304 62698 108356 62704
rect 109328 62490 109356 65484
rect 109316 62484 109368 62490
rect 109316 62426 109368 62432
rect 108304 62348 108356 62354
rect 108304 62290 108356 62296
rect 107384 61396 107436 61402
rect 107384 61338 107436 61344
rect 108120 3868 108172 3874
rect 108120 3810 108172 3816
rect 107016 3392 107068 3398
rect 107016 3334 107068 3340
rect 108132 480 108160 3810
rect 108316 3806 108344 62290
rect 110248 61538 110276 65484
rect 111260 62558 111288 65484
rect 112180 62898 112208 65484
rect 112168 62892 112220 62898
rect 112168 62834 112220 62840
rect 113088 62892 113140 62898
rect 113088 62834 113140 62840
rect 111248 62552 111300 62558
rect 111248 62494 111300 62500
rect 112444 62484 112496 62490
rect 112444 62426 112496 62432
rect 110236 61532 110288 61538
rect 110236 61474 110288 61480
rect 111708 61396 111760 61402
rect 111708 61338 111760 61344
rect 111720 6914 111748 61338
rect 111628 6886 111748 6914
rect 109316 3868 109368 3874
rect 109316 3810 109368 3816
rect 108304 3800 108356 3806
rect 108304 3742 108356 3748
rect 109328 480 109356 3810
rect 110512 3664 110564 3670
rect 110512 3606 110564 3612
rect 110524 480 110552 3606
rect 111628 480 111656 6886
rect 112456 3194 112484 62426
rect 113100 6914 113128 62834
rect 113192 61470 113220 65484
rect 113824 62416 113876 62422
rect 113824 62358 113876 62364
rect 113180 61464 113232 61470
rect 113180 61406 113232 61412
rect 112824 6886 113128 6914
rect 112444 3188 112496 3194
rect 112444 3130 112496 3136
rect 112824 480 112852 6886
rect 113836 4010 113864 62358
rect 114112 62286 114140 65484
rect 114100 62280 114152 62286
rect 114100 62222 114152 62228
rect 115124 62218 115152 65484
rect 115848 63436 115900 63442
rect 115848 63378 115900 63384
rect 115112 62212 115164 62218
rect 115112 62154 115164 62160
rect 113916 62144 113968 62150
rect 113916 62086 113968 62092
rect 113824 4004 113876 4010
rect 113824 3946 113876 3952
rect 113928 3602 113956 62086
rect 114008 3800 114060 3806
rect 114008 3742 114060 3748
rect 113916 3596 113968 3602
rect 113916 3538 113968 3544
rect 114020 480 114048 3742
rect 115860 3602 115888 63378
rect 116044 61606 116072 65484
rect 117056 63510 117084 65484
rect 117044 63504 117096 63510
rect 117044 63446 117096 63452
rect 117228 62756 117280 62762
rect 117228 62698 117280 62704
rect 116584 62552 116636 62558
rect 116584 62494 116636 62500
rect 116032 61600 116084 61606
rect 116032 61542 116084 61548
rect 116596 3874 116624 62494
rect 116584 3868 116636 3874
rect 116584 3810 116636 3816
rect 117240 3602 117268 62698
rect 117976 62354 118004 65484
rect 117964 62348 118016 62354
rect 117964 62290 118016 62296
rect 118988 61878 119016 65484
rect 119804 63504 119856 63510
rect 119804 63446 119856 63452
rect 118976 61872 119028 61878
rect 118976 61814 119028 61820
rect 119816 55214 119844 63446
rect 119908 63034 119936 65484
rect 119896 63028 119948 63034
rect 119896 62970 119948 62976
rect 119988 63028 120040 63034
rect 119988 62970 120040 62976
rect 119816 55186 119936 55214
rect 119908 16574 119936 55186
rect 119816 16546 119936 16574
rect 117596 3868 117648 3874
rect 117596 3810 117648 3816
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 115216 480 115244 3538
rect 116412 480 116440 3538
rect 117608 480 117636 3810
rect 119816 3602 119844 16546
rect 120000 6914 120028 62970
rect 120724 62280 120776 62286
rect 120724 62222 120776 62228
rect 119908 6886 120028 6914
rect 118792 3596 118844 3602
rect 118792 3538 118844 3544
rect 119804 3596 119856 3602
rect 119804 3538 119856 3544
rect 118804 480 118832 3538
rect 119908 480 119936 6886
rect 120736 4078 120764 62222
rect 120920 62150 120948 65484
rect 120908 62144 120960 62150
rect 120908 62086 120960 62092
rect 121840 61946 121868 65484
rect 122748 62688 122800 62694
rect 122748 62630 122800 62636
rect 121828 61940 121880 61946
rect 121828 61882 121880 61888
rect 120724 4072 120776 4078
rect 120724 4014 120776 4020
rect 122760 3602 122788 62630
rect 122852 62626 122880 65484
rect 123772 63170 123800 65484
rect 123760 63164 123812 63170
rect 123760 63106 123812 63112
rect 124128 63164 124180 63170
rect 124128 63106 124180 63112
rect 122840 62620 122892 62626
rect 122840 62562 122892 62568
rect 123484 62348 123536 62354
rect 123484 62290 123536 62296
rect 123496 6914 123524 62290
rect 123404 6886 123524 6914
rect 123404 4146 123432 6886
rect 123392 4140 123444 4146
rect 123392 4082 123444 4088
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 121092 3392 121144 3398
rect 121092 3334 121144 3340
rect 121104 480 121132 3334
rect 122300 480 122328 3538
rect 124140 3330 124168 63106
rect 124784 6254 124812 65484
rect 125704 62966 125732 65484
rect 125692 62960 125744 62966
rect 125692 62902 125744 62908
rect 125508 62620 125560 62626
rect 125508 62562 125560 62568
rect 124772 6248 124824 6254
rect 124772 6190 124824 6196
rect 125520 3602 125548 62562
rect 126716 62422 126744 65484
rect 126704 62416 126756 62422
rect 126704 62358 126756 62364
rect 127636 62014 127664 65484
rect 128648 62490 128676 65484
rect 129568 63238 129596 65484
rect 129556 63232 129608 63238
rect 129556 63174 129608 63180
rect 129004 62960 129056 62966
rect 129004 62902 129056 62908
rect 128636 62484 128688 62490
rect 128636 62426 128688 62432
rect 127624 62008 127676 62014
rect 127624 61950 127676 61956
rect 126888 61464 126940 61470
rect 126888 61406 126940 61412
rect 126900 3602 126928 61406
rect 128360 4888 128412 4894
rect 128360 4830 128412 4836
rect 128176 4004 128228 4010
rect 128176 3946 128228 3952
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 125508 3596 125560 3602
rect 125508 3538 125560 3544
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 126888 3596 126940 3602
rect 126888 3538 126940 3544
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 123484 3324 123536 3330
rect 123484 3266 123536 3272
rect 124128 3324 124180 3330
rect 124128 3266 124180 3272
rect 123496 480 123524 3266
rect 124692 480 124720 3538
rect 125888 480 125916 3538
rect 126992 480 127020 3538
rect 128188 480 128216 3946
rect 128372 3942 128400 4830
rect 128360 3936 128412 3942
rect 128360 3878 128412 3884
rect 129016 3738 129044 62902
rect 130580 61674 130608 65484
rect 131500 63102 131528 65484
rect 131488 63096 131540 63102
rect 131488 63038 131540 63044
rect 132512 62286 132540 65484
rect 132500 62280 132552 62286
rect 132500 62222 132552 62228
rect 133144 62212 133196 62218
rect 133144 62154 133196 62160
rect 130568 61668 130620 61674
rect 130568 61610 130620 61616
rect 131028 61532 131080 61538
rect 131028 61474 131080 61480
rect 130384 61328 130436 61334
rect 130384 61270 130436 61276
rect 129372 6248 129424 6254
rect 129372 6190 129424 6196
rect 129004 3732 129056 3738
rect 129004 3674 129056 3680
rect 129384 480 129412 6190
rect 130396 3602 130424 61270
rect 131040 3602 131068 61474
rect 132960 3732 133012 3738
rect 132960 3674 133012 3680
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 130568 3596 130620 3602
rect 130568 3538 130620 3544
rect 131028 3596 131080 3602
rect 131028 3538 131080 3544
rect 130580 480 130608 3538
rect 131764 3324 131816 3330
rect 131764 3266 131816 3272
rect 131776 480 131804 3266
rect 132972 480 133000 3674
rect 133156 3534 133184 62154
rect 133432 61810 133460 65484
rect 134444 63306 134472 65484
rect 134432 63300 134484 63306
rect 134432 63242 134484 63248
rect 134524 63232 134576 63238
rect 134524 63174 134576 63180
rect 133420 61804 133472 61810
rect 133420 61746 133472 61752
rect 133236 61600 133288 61606
rect 133236 61542 133288 61548
rect 133144 3528 133196 3534
rect 133144 3470 133196 3476
rect 133248 3330 133276 61542
rect 134536 3670 134564 63174
rect 135364 62354 135392 65484
rect 135904 62416 135956 62422
rect 135904 62358 135956 62364
rect 135352 62348 135404 62354
rect 135352 62290 135404 62296
rect 134616 62144 134668 62150
rect 134616 62086 134668 62092
rect 134628 6186 134656 62086
rect 134616 6180 134668 6186
rect 134616 6122 134668 6128
rect 135916 3806 135944 62358
rect 136376 62150 136404 65484
rect 137296 62830 137324 65484
rect 138308 62966 138336 65484
rect 138664 63300 138716 63306
rect 138664 63242 138716 63248
rect 138296 62960 138348 62966
rect 138296 62902 138348 62908
rect 137284 62824 137336 62830
rect 137284 62766 137336 62772
rect 137284 62484 137336 62490
rect 137284 62426 137336 62432
rect 136364 62144 136416 62150
rect 136364 62086 136416 62092
rect 137296 3874 137324 62426
rect 137376 62144 137428 62150
rect 137376 62086 137428 62092
rect 137284 3868 137336 3874
rect 137284 3810 137336 3816
rect 135904 3800 135956 3806
rect 135904 3742 135956 3748
rect 134524 3664 134576 3670
rect 134524 3606 134576 3612
rect 134156 3596 134208 3602
rect 134156 3538 134208 3544
rect 133236 3324 133288 3330
rect 133236 3266 133288 3272
rect 134168 480 134196 3538
rect 137388 3534 137416 62086
rect 137376 3528 137428 3534
rect 137376 3470 137428 3476
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135272 480 135300 3402
rect 138676 3398 138704 63242
rect 139228 62150 139256 65484
rect 140240 63374 140268 65484
rect 140228 63368 140280 63374
rect 140228 63310 140280 63316
rect 139308 62824 139360 62830
rect 139308 62766 139360 62772
rect 139216 62144 139268 62150
rect 139216 62086 139268 62092
rect 138664 3392 138716 3398
rect 138664 3334 138716 3340
rect 139320 3330 139348 62766
rect 141160 62218 141188 65484
rect 142068 63096 142120 63102
rect 142068 63038 142120 63044
rect 141148 62212 141200 62218
rect 141148 62154 141200 62160
rect 141424 61940 141476 61946
rect 141424 61882 141476 61888
rect 140688 61736 140740 61742
rect 140688 61678 140740 61684
rect 139400 4820 139452 4826
rect 139400 4762 139452 4768
rect 138848 3324 138900 3330
rect 138848 3266 138900 3272
rect 139308 3324 139360 3330
rect 139308 3266 139360 3272
rect 136456 3256 136508 3262
rect 136456 3198 136508 3204
rect 136468 480 136496 3198
rect 137652 2848 137704 2854
rect 137652 2790 137704 2796
rect 137664 480 137692 2790
rect 138860 480 138888 3266
rect 139412 2854 139440 4762
rect 140700 3534 140728 61678
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 139400 2848 139452 2854
rect 139400 2790 139452 2796
rect 140056 480 140084 3470
rect 141240 3460 141292 3466
rect 141240 3402 141292 3408
rect 141252 480 141280 3402
rect 141436 3262 141464 61882
rect 142080 3466 142108 63038
rect 142172 4894 142200 65484
rect 143092 62558 143120 65484
rect 144104 63238 144132 65484
rect 145024 64874 145052 65484
rect 144932 64846 145052 64874
rect 144932 63322 144960 64846
rect 144656 63294 144960 63322
rect 144092 63232 144144 63238
rect 144092 63174 144144 63180
rect 143448 62960 143500 62966
rect 143448 62902 143500 62908
rect 143080 62552 143132 62558
rect 143080 62494 143132 62500
rect 142160 4888 142212 4894
rect 142160 4830 142212 4836
rect 143460 3466 143488 62902
rect 144656 61402 144684 63294
rect 144828 63232 144880 63238
rect 144828 63174 144880 63180
rect 144644 61396 144696 61402
rect 144644 61338 144696 61344
rect 144736 61396 144788 61402
rect 144736 61338 144788 61344
rect 144748 16574 144776 61338
rect 144656 16546 144776 16574
rect 144656 3466 144684 16546
rect 144840 6914 144868 63174
rect 146036 62898 146064 65484
rect 146956 64874 146984 65484
rect 146864 64846 146984 64874
rect 146024 62892 146076 62898
rect 146024 62834 146076 62840
rect 146864 62422 146892 64846
rect 147968 63442 147996 65484
rect 147956 63436 148008 63442
rect 147956 63378 148008 63384
rect 148888 62762 148916 65484
rect 148968 63368 149020 63374
rect 148968 63310 149020 63316
rect 148876 62756 148928 62762
rect 148876 62698 148928 62704
rect 146944 62552 146996 62558
rect 146944 62494 146996 62500
rect 146852 62416 146904 62422
rect 146852 62358 146904 62364
rect 144748 6886 144868 6914
rect 142068 3460 142120 3466
rect 142068 3402 142120 3408
rect 142436 3460 142488 3466
rect 142436 3402 142488 3408
rect 143448 3460 143500 3466
rect 143448 3402 143500 3408
rect 143540 3460 143592 3466
rect 143540 3402 143592 3408
rect 144644 3460 144696 3466
rect 144644 3402 144696 3408
rect 141424 3256 141476 3262
rect 141424 3198 141476 3204
rect 142448 480 142476 3402
rect 143552 480 143580 3402
rect 144748 480 144776 6886
rect 146956 4010 146984 62494
rect 147588 61804 147640 61810
rect 147588 61746 147640 61752
rect 146944 4004 146996 4010
rect 146944 3946 146996 3952
rect 147600 3466 147628 61746
rect 148980 3466 149008 63310
rect 149900 62490 149928 65484
rect 150820 63510 150848 65484
rect 150808 63504 150860 63510
rect 150808 63446 150860 63452
rect 151832 63034 151860 65484
rect 152752 63306 152780 65484
rect 153016 63436 153068 63442
rect 153016 63378 153068 63384
rect 152740 63300 152792 63306
rect 152740 63242 152792 63248
rect 151820 63028 151872 63034
rect 151820 62970 151872 62976
rect 150348 62892 150400 62898
rect 150348 62834 150400 62840
rect 149888 62484 149940 62490
rect 149888 62426 149940 62432
rect 150360 3466 150388 62834
rect 151084 62008 151136 62014
rect 151084 61950 151136 61956
rect 151096 3738 151124 61950
rect 151728 61872 151780 61878
rect 151728 61814 151780 61820
rect 151084 3732 151136 3738
rect 151084 3674 151136 3680
rect 151740 3466 151768 61814
rect 153028 16574 153056 63378
rect 153108 63028 153160 63034
rect 153108 62970 153160 62976
rect 152936 16546 153056 16574
rect 147128 3460 147180 3466
rect 147128 3402 147180 3408
rect 147588 3460 147640 3466
rect 147588 3402 147640 3408
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148968 3460 149020 3466
rect 148968 3402 149020 3408
rect 149520 3460 149572 3466
rect 149520 3402 149572 3408
rect 150348 3460 150400 3466
rect 150348 3402 150400 3408
rect 150624 3460 150676 3466
rect 150624 3402 150676 3408
rect 151728 3460 151780 3466
rect 151728 3402 151780 3408
rect 145932 3392 145984 3398
rect 145932 3334 145984 3340
rect 145944 480 145972 3334
rect 147140 480 147168 3402
rect 148336 480 148364 3402
rect 149532 480 149560 3402
rect 150636 480 150664 3402
rect 152936 3058 152964 16546
rect 153120 6914 153148 62970
rect 153764 62694 153792 65484
rect 154488 63300 154540 63306
rect 154488 63242 154540 63248
rect 153752 62688 153804 62694
rect 153752 62630 153804 62636
rect 154500 6914 154528 63242
rect 154684 63170 154712 65484
rect 154672 63164 154724 63170
rect 154672 63106 154724 63112
rect 155696 62626 155724 65484
rect 156616 64874 156644 65484
rect 156524 64846 156644 64874
rect 155868 63164 155920 63170
rect 155868 63106 155920 63112
rect 155684 62620 155736 62626
rect 155684 62562 155736 62568
rect 155224 61260 155276 61266
rect 155224 61202 155276 61208
rect 153028 6886 153148 6914
rect 154224 6886 154528 6914
rect 151820 3052 151872 3058
rect 151820 2994 151872 3000
rect 152924 3052 152976 3058
rect 152924 2994 152976 3000
rect 151832 480 151860 2994
rect 153028 480 153056 6886
rect 154224 480 154252 6886
rect 155236 3602 155264 61202
rect 155224 3596 155276 3602
rect 155224 3538 155276 3544
rect 155880 3534 155908 63106
rect 156524 61470 156552 64846
rect 157248 63504 157300 63510
rect 157248 63446 157300 63452
rect 156604 62416 156656 62422
rect 156604 62358 156656 62364
rect 156512 61464 156564 61470
rect 156512 61406 156564 61412
rect 156616 3670 156644 62358
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 157260 3534 157288 63446
rect 157628 61334 157656 65484
rect 158548 62558 158576 65484
rect 158628 62688 158680 62694
rect 158628 62630 158680 62636
rect 158536 62552 158588 62558
rect 158536 62494 158588 62500
rect 157616 61328 157668 61334
rect 157616 61270 157668 61276
rect 158640 3534 158668 62630
rect 159560 6254 159588 65484
rect 160008 62620 160060 62626
rect 160008 62562 160060 62568
rect 159548 6248 159600 6254
rect 159548 6190 159600 6196
rect 160020 3534 160048 62562
rect 160480 61538 160508 65484
rect 161388 62484 161440 62490
rect 161388 62426 161440 62432
rect 160744 62348 160796 62354
rect 160744 62290 160796 62296
rect 160468 61532 160520 61538
rect 160468 61474 160520 61480
rect 155408 3528 155460 3534
rect 155408 3470 155460 3476
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 155420 480 155448 3470
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3470
rect 160756 3398 160784 62290
rect 161296 4140 161348 4146
rect 161296 4082 161348 4088
rect 160744 3392 160796 3398
rect 160744 3334 160796 3340
rect 161308 480 161336 4082
rect 161400 3534 161428 62426
rect 161492 61606 161520 65484
rect 162412 62014 162440 65484
rect 162768 62756 162820 62762
rect 162768 62698 162820 62704
rect 162400 62008 162452 62014
rect 162400 61950 162452 61956
rect 161480 61600 161532 61606
rect 161480 61542 161532 61548
rect 162124 61464 162176 61470
rect 162124 61406 162176 61412
rect 162136 4146 162164 61406
rect 162780 6914 162808 62698
rect 163424 61266 163452 65484
rect 164148 62552 164200 62558
rect 164148 62494 164200 62500
rect 163412 61260 163464 61266
rect 163412 61202 163464 61208
rect 162504 6886 162808 6914
rect 162124 4140 162176 4146
rect 162124 4082 162176 4088
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 162504 480 162532 6886
rect 164160 3330 164188 62494
rect 164344 62422 164372 65484
rect 164332 62416 164384 62422
rect 164332 62358 164384 62364
rect 165356 61946 165384 65484
rect 165344 61940 165396 61946
rect 165344 61882 165396 61888
rect 165528 61532 165580 61538
rect 165528 61474 165580 61480
rect 165540 3534 165568 61474
rect 166276 4826 166304 65484
rect 167288 62830 167316 65484
rect 167276 62824 167328 62830
rect 167276 62766 167328 62772
rect 166908 62416 166960 62422
rect 166908 62358 166960 62364
rect 166264 4820 166316 4826
rect 166264 4762 166316 4768
rect 166920 3534 166948 62358
rect 168208 61742 168236 65484
rect 169220 63102 169248 65484
rect 169208 63096 169260 63102
rect 169208 63038 169260 63044
rect 169668 63096 169720 63102
rect 169668 63038 169720 63044
rect 168288 62824 168340 62830
rect 168288 62766 168340 62772
rect 168196 61736 168248 61742
rect 168196 61678 168248 61684
rect 168300 3534 168328 62766
rect 169680 6914 169708 63038
rect 170140 62966 170168 65484
rect 170128 62960 170180 62966
rect 170128 62902 170180 62908
rect 171048 62960 171100 62966
rect 171048 62902 171100 62908
rect 171060 6914 171088 62902
rect 171152 61402 171180 65484
rect 172072 63238 172100 65484
rect 172060 63232 172112 63238
rect 172060 63174 172112 63180
rect 173084 62354 173112 65484
rect 173072 62348 173124 62354
rect 173072 62290 173124 62296
rect 173808 62348 173860 62354
rect 173808 62290 173860 62296
rect 171140 61396 171192 61402
rect 171140 61338 171192 61344
rect 173164 61396 173216 61402
rect 173164 61338 173216 61344
rect 169588 6886 169708 6914
rect 170784 6886 171088 6914
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 165528 3528 165580 3534
rect 165528 3470 165580 3476
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 168288 3528 168340 3534
rect 168288 3470 168340 3476
rect 163688 3324 163740 3330
rect 163688 3266 163740 3272
rect 164148 3324 164200 3330
rect 164148 3266 164200 3272
rect 163700 480 163728 3266
rect 164896 480 164924 3470
rect 166092 480 166120 3470
rect 167196 480 167224 3470
rect 168380 3120 168432 3126
rect 168380 3062 168432 3068
rect 168392 480 168420 3062
rect 169588 480 169616 6886
rect 169760 6180 169812 6186
rect 169760 6122 169812 6128
rect 169772 3126 169800 6122
rect 169760 3120 169812 3126
rect 169760 3062 169812 3068
rect 170784 480 170812 6886
rect 173176 3670 173204 61338
rect 171968 3664 172020 3670
rect 171968 3606 172020 3612
rect 173164 3664 173216 3670
rect 173164 3606 173216 3612
rect 171980 480 172008 3606
rect 173820 3534 173848 62290
rect 174004 61810 174032 65484
rect 175016 63374 175044 65484
rect 175004 63368 175056 63374
rect 175004 63310 175056 63316
rect 175188 63232 175240 63238
rect 175188 63174 175240 63180
rect 173992 61804 174044 61810
rect 173992 61746 174044 61752
rect 175200 3534 175228 63174
rect 175936 62898 175964 65484
rect 175924 62892 175976 62898
rect 175924 62834 175976 62840
rect 176568 62280 176620 62286
rect 176568 62222 176620 62228
rect 176580 3534 176608 62222
rect 176948 61878 176976 65484
rect 177868 63442 177896 65484
rect 177856 63436 177908 63442
rect 177856 63378 177908 63384
rect 177948 63368 178000 63374
rect 177948 63310 178000 63316
rect 177856 62892 177908 62898
rect 177856 62834 177908 62840
rect 176936 61872 176988 61878
rect 176936 61814 176988 61820
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 173176 480 173204 3470
rect 174280 480 174308 3470
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 62834
rect 177960 3534 177988 63310
rect 178880 63034 178908 65484
rect 179800 63306 179828 65484
rect 179788 63300 179840 63306
rect 179788 63242 179840 63248
rect 180708 63300 180760 63306
rect 180708 63242 180760 63248
rect 178868 63028 178920 63034
rect 178868 62970 178920 62976
rect 179328 63028 179380 63034
rect 179328 62970 179380 62976
rect 179340 6914 179368 62970
rect 179064 6886 179368 6914
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179064 480 179092 6886
rect 180720 3534 180748 63242
rect 180812 63170 180840 65484
rect 181732 63510 181760 65484
rect 181720 63504 181772 63510
rect 181720 63446 181772 63452
rect 180800 63164 180852 63170
rect 180800 63106 180852 63112
rect 182088 63164 182140 63170
rect 182088 63106 182140 63112
rect 182100 3534 182128 63106
rect 182744 62694 182772 65484
rect 183468 63504 183520 63510
rect 183468 63446 183520 63452
rect 182732 62688 182784 62694
rect 182732 62630 182784 62636
rect 183480 3534 183508 63446
rect 183664 62626 183692 65484
rect 183652 62620 183704 62626
rect 183652 62562 183704 62568
rect 184676 62490 184704 65484
rect 184848 62620 184900 62626
rect 184848 62562 184900 62568
rect 184664 62484 184716 62490
rect 184664 62426 184716 62432
rect 184860 3534 184888 62562
rect 185596 61470 185624 65484
rect 186228 63436 186280 63442
rect 186228 63378 186280 63384
rect 185584 61464 185636 61470
rect 185584 61406 185636 61412
rect 186240 6914 186268 63378
rect 186608 62762 186636 65484
rect 186596 62756 186648 62762
rect 186596 62698 186648 62704
rect 187528 62558 187556 65484
rect 187516 62552 187568 62558
rect 187516 62494 187568 62500
rect 187608 62552 187660 62558
rect 187608 62494 187660 62500
rect 187620 6914 187648 62494
rect 188344 62212 188396 62218
rect 188344 62154 188396 62160
rect 186148 6886 186268 6914
rect 187344 6886 187648 6914
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182560 480 182588 3470
rect 183756 480 183784 3470
rect 184940 3324 184992 3330
rect 184940 3266 184992 3272
rect 184952 480 184980 3266
rect 186148 480 186176 6886
rect 187344 480 187372 6886
rect 188356 3330 188384 62154
rect 188540 61538 188568 65484
rect 188988 62756 189040 62762
rect 188988 62698 189040 62704
rect 188528 61532 188580 61538
rect 188528 61474 188580 61480
rect 189000 3534 189028 62698
rect 189460 62422 189488 65484
rect 190472 62830 190500 65484
rect 190460 62824 190512 62830
rect 190460 62766 190512 62772
rect 190368 62688 190420 62694
rect 190368 62630 190420 62636
rect 189448 62416 189500 62422
rect 189448 62358 189500 62364
rect 190380 3534 190408 62630
rect 191392 6186 191420 65484
rect 192404 63102 192432 65484
rect 192392 63096 192444 63102
rect 192392 63038 192444 63044
rect 193324 62966 193352 65484
rect 193312 62960 193364 62966
rect 193312 62902 193364 62908
rect 191748 62824 191800 62830
rect 191748 62766 191800 62772
rect 191380 6180 191432 6186
rect 191380 6122 191432 6128
rect 191760 3534 191788 62766
rect 193128 62416 193180 62422
rect 193128 62358 193180 62364
rect 193140 3534 193168 62358
rect 194336 61402 194364 65484
rect 194416 63096 194468 63102
rect 194416 63038 194468 63044
rect 194324 61396 194376 61402
rect 194324 61338 194376 61344
rect 194428 16574 194456 63038
rect 194508 62960 194560 62966
rect 194508 62902 194560 62908
rect 194336 16546 194456 16574
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 189724 3528 189776 3534
rect 189724 3470 189776 3476
rect 190368 3528 190420 3534
rect 190368 3470 190420 3476
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 188344 3324 188396 3330
rect 188344 3266 188396 3272
rect 188540 480 188568 3470
rect 189736 480 189764 3470
rect 190840 480 190868 3470
rect 192036 480 192064 3470
rect 194336 3194 194364 16546
rect 194520 6914 194548 62902
rect 195256 62354 195284 65484
rect 196268 63238 196296 65484
rect 196256 63232 196308 63238
rect 196256 63174 196308 63180
rect 195888 62484 195940 62490
rect 195888 62426 195940 62432
rect 195244 62348 195296 62354
rect 195244 62290 195296 62296
rect 195900 6914 195928 62426
rect 197188 62286 197216 65484
rect 198200 63374 198228 65484
rect 198188 63368 198240 63374
rect 198188 63310 198240 63316
rect 198648 63368 198700 63374
rect 198648 63310 198700 63316
rect 197268 63232 197320 63238
rect 197268 63174 197320 63180
rect 197176 62280 197228 62286
rect 197176 62222 197228 62228
rect 194428 6886 194548 6914
rect 195624 6886 195928 6914
rect 193220 3188 193272 3194
rect 193220 3130 193272 3136
rect 194324 3188 194376 3194
rect 194324 3130 194376 3136
rect 193232 480 193260 3130
rect 194428 480 194456 6886
rect 195624 480 195652 6886
rect 197280 3058 197308 63174
rect 198660 3534 198688 63310
rect 199120 62898 199148 65484
rect 200132 63034 200160 65484
rect 201052 63306 201080 65484
rect 201040 63300 201092 63306
rect 201040 63242 201092 63248
rect 202064 63170 202092 65484
rect 202984 63510 203012 65484
rect 202972 63504 203024 63510
rect 202972 63446 203024 63452
rect 202052 63164 202104 63170
rect 202052 63106 202104 63112
rect 200120 63028 200172 63034
rect 200120 62970 200172 62976
rect 199108 62892 199160 62898
rect 199108 62834 199160 62840
rect 202696 62892 202748 62898
rect 202696 62834 202748 62840
rect 200028 62348 200080 62354
rect 200028 62290 200080 62296
rect 200040 3534 200068 62290
rect 201408 62280 201460 62286
rect 201408 62222 201460 62228
rect 201420 3534 201448 62222
rect 197912 3528 197964 3534
rect 197912 3470 197964 3476
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 200304 3528 200356 3534
rect 200304 3470 200356 3476
rect 201408 3528 201460 3534
rect 201408 3470 201460 3476
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 196808 3052 196860 3058
rect 196808 2994 196860 3000
rect 197268 3052 197320 3058
rect 197268 2994 197320 3000
rect 196820 480 196848 2994
rect 197924 480 197952 3470
rect 199120 480 199148 3470
rect 200316 480 200344 3470
rect 201512 480 201540 3470
rect 202708 480 202736 62834
rect 203996 62626 204024 65484
rect 204168 63300 204220 63306
rect 204168 63242 204220 63248
rect 203984 62620 204036 62626
rect 203984 62562 204036 62568
rect 202788 62144 202840 62150
rect 202788 62086 202840 62092
rect 202800 3534 202828 62086
rect 204180 6914 204208 63242
rect 204916 62218 204944 65484
rect 205928 63442 205956 65484
rect 205916 63436 205968 63442
rect 205916 63378 205968 63384
rect 205548 63164 205600 63170
rect 205548 63106 205600 63112
rect 204904 62212 204956 62218
rect 204904 62154 204956 62160
rect 203904 6886 204208 6914
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 203904 480 203932 6886
rect 205560 3534 205588 63106
rect 206848 62558 206876 65484
rect 206928 63028 206980 63034
rect 206928 62970 206980 62976
rect 206836 62552 206888 62558
rect 206836 62494 206888 62500
rect 206940 3534 206968 62970
rect 207860 62762 207888 65484
rect 207848 62756 207900 62762
rect 207848 62698 207900 62704
rect 208308 62756 208360 62762
rect 208308 62698 208360 62704
rect 208320 3534 208348 62698
rect 208780 62694 208808 65484
rect 209688 63504 209740 63510
rect 209688 63446 209740 63452
rect 208768 62688 208820 62694
rect 208768 62630 208820 62636
rect 209700 3534 209728 63446
rect 209792 62830 209820 65484
rect 209780 62824 209832 62830
rect 209780 62766 209832 62772
rect 210712 62422 210740 65484
rect 211068 63436 211120 63442
rect 211068 63378 211120 63384
rect 210976 62824 211028 62830
rect 210976 62766 211028 62772
rect 210700 62416 210752 62422
rect 210700 62358 210752 62364
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207400 480 207428 3470
rect 208596 480 208624 3470
rect 209792 480 209820 3470
rect 210988 480 211016 62766
rect 211080 3534 211108 63378
rect 211724 63102 211752 65484
rect 211712 63096 211764 63102
rect 211712 63038 211764 63044
rect 212448 63096 212500 63102
rect 212448 63038 212500 63044
rect 212460 6914 212488 63038
rect 212644 62966 212672 65484
rect 212632 62960 212684 62966
rect 212632 62902 212684 62908
rect 213656 62490 213684 65484
rect 214576 63238 214604 65484
rect 215588 63374 215616 65484
rect 215576 63368 215628 63374
rect 215576 63310 215628 63316
rect 214564 63232 214616 63238
rect 214564 63174 214616 63180
rect 215208 63232 215260 63238
rect 215208 63174 215260 63180
rect 213828 62960 213880 62966
rect 213828 62902 213880 62908
rect 213644 62484 213696 62490
rect 213644 62426 213696 62432
rect 212184 6886 212488 6914
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 212184 480 212212 6886
rect 213840 3534 213868 62902
rect 215220 3534 215248 63174
rect 216508 62354 216536 65484
rect 216588 62552 216640 62558
rect 216588 62494 216640 62500
rect 216496 62348 216548 62354
rect 216496 62290 216548 62296
rect 216600 3534 216628 62494
rect 217520 62286 217548 65484
rect 217968 62688 218020 62694
rect 217968 62630 218020 62636
rect 217508 62280 217560 62286
rect 217508 62222 217560 62228
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 213380 480 213408 3470
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 217980 3194 218008 62630
rect 218440 62150 218468 65484
rect 219256 63368 219308 63374
rect 219256 63310 219308 63316
rect 218428 62144 218480 62150
rect 218428 62086 218480 62092
rect 219268 16574 219296 63310
rect 219452 62898 219480 65484
rect 220372 63306 220400 65484
rect 220360 63300 220412 63306
rect 220360 63242 220412 63248
rect 221384 63170 221412 65484
rect 221372 63164 221424 63170
rect 221372 63106 221424 63112
rect 222108 63164 222160 63170
rect 222108 63106 222160 63112
rect 219440 62892 219492 62898
rect 219440 62834 219492 62840
rect 220728 62892 220780 62898
rect 220728 62834 220780 62840
rect 219348 62620 219400 62626
rect 219348 62562 219400 62568
rect 219176 16546 219296 16574
rect 219176 3534 219204 16546
rect 219360 6914 219388 62562
rect 220740 6914 220768 62834
rect 219268 6886 219388 6914
rect 220464 6886 220768 6914
rect 218060 3528 218112 3534
rect 218060 3470 218112 3476
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 216864 3188 216916 3194
rect 216864 3130 216916 3136
rect 217968 3188 218020 3194
rect 217968 3130 218020 3136
rect 216876 480 216904 3130
rect 218072 480 218100 3470
rect 219268 480 219296 6886
rect 220464 480 220492 6886
rect 222120 3126 222148 63106
rect 222304 63034 222332 65484
rect 222292 63028 222344 63034
rect 222292 62970 222344 62976
rect 223316 62762 223344 65484
rect 224236 63510 224264 65484
rect 224224 63504 224276 63510
rect 224224 63446 224276 63452
rect 225248 63442 225276 65484
rect 225236 63436 225288 63442
rect 225236 63378 225288 63384
rect 223488 63300 223540 63306
rect 223488 63242 223540 63248
rect 223304 62756 223356 62762
rect 223304 62698 223356 62704
rect 223500 3534 223528 63242
rect 224868 63028 224920 63034
rect 224868 62970 224920 62976
rect 224880 3534 224908 62970
rect 226168 62830 226196 65484
rect 226248 63436 226300 63442
rect 226248 63378 226300 63384
rect 226156 62824 226208 62830
rect 226156 62766 226208 62772
rect 226260 3534 226288 63378
rect 227180 63102 227208 65484
rect 227168 63096 227220 63102
rect 227168 63038 227220 63044
rect 227628 63096 227680 63102
rect 227628 63038 227680 63044
rect 227536 62824 227588 62830
rect 227536 62766 227588 62772
rect 227548 16574 227576 62766
rect 227456 16546 227576 16574
rect 227456 3534 227484 16546
rect 227640 6914 227668 63038
rect 228100 62966 228128 65484
rect 229008 63504 229060 63510
rect 229008 63446 229060 63452
rect 228088 62960 228140 62966
rect 228088 62902 228140 62908
rect 229020 6914 229048 63446
rect 229112 63238 229140 65484
rect 229100 63232 229152 63238
rect 229100 63174 229152 63180
rect 230032 62558 230060 65484
rect 230388 62960 230440 62966
rect 230388 62902 230440 62908
rect 230020 62552 230072 62558
rect 230020 62494 230072 62500
rect 227548 6886 227668 6914
rect 228744 6886 229048 6914
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 225144 3528 225196 3534
rect 225144 3470 225196 3476
rect 226248 3528 226300 3534
rect 226248 3470 226300 3476
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 227444 3528 227496 3534
rect 227444 3470 227496 3476
rect 221556 3120 221608 3126
rect 221556 3062 221608 3068
rect 222108 3120 222160 3126
rect 222108 3062 222160 3068
rect 221568 480 221596 3062
rect 222764 480 222792 3470
rect 223960 480 223988 3470
rect 225156 480 225184 3470
rect 226352 480 226380 3470
rect 227548 480 227576 6886
rect 228744 480 228772 6886
rect 230400 3330 230428 62902
rect 231044 62694 231072 65484
rect 231964 63374 231992 65484
rect 231952 63368 232004 63374
rect 231952 63310 232004 63316
rect 231768 63232 231820 63238
rect 231768 63174 231820 63180
rect 231032 62688 231084 62694
rect 231032 62630 231084 62636
rect 231780 3534 231808 63174
rect 232976 62626 233004 65484
rect 233148 63368 233200 63374
rect 233148 63310 233200 63316
rect 232964 62620 233016 62626
rect 232964 62562 233016 62568
rect 233160 3534 233188 63310
rect 233896 62898 233924 65484
rect 234908 63170 234936 65484
rect 235828 63306 235856 65484
rect 235816 63300 235868 63306
rect 235816 63242 235868 63248
rect 235908 63300 235960 63306
rect 235908 63242 235960 63248
rect 234896 63164 234948 63170
rect 234896 63106 234948 63112
rect 233884 62892 233936 62898
rect 233884 62834 233936 62840
rect 234528 62892 234580 62898
rect 234528 62834 234580 62840
rect 234540 3534 234568 62834
rect 235816 62756 235868 62762
rect 235816 62698 235868 62704
rect 235828 16574 235856 62698
rect 235736 16546 235856 16574
rect 235736 3534 235764 16546
rect 235920 6914 235948 63242
rect 236840 63034 236868 65484
rect 237760 63442 237788 65484
rect 237748 63436 237800 63442
rect 237748 63378 237800 63384
rect 237288 63164 237340 63170
rect 237288 63106 237340 63112
rect 236828 63028 236880 63034
rect 236828 62970 236880 62976
rect 237300 6914 237328 63106
rect 238668 63028 238720 63034
rect 238668 62970 238720 62976
rect 235828 6886 235948 6914
rect 237024 6886 237328 6914
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 235724 3528 235776 3534
rect 235724 3470 235776 3476
rect 229836 3324 229888 3330
rect 229836 3266 229888 3272
rect 230388 3324 230440 3330
rect 230388 3266 230440 3272
rect 229848 480 229876 3266
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235828 480 235856 6886
rect 237024 480 237052 6886
rect 238680 3330 238708 62970
rect 238772 62830 238800 65484
rect 239692 63102 239720 65484
rect 240704 63510 240732 65484
rect 240692 63504 240744 63510
rect 240692 63446 240744 63452
rect 240784 63436 240836 63442
rect 240784 63378 240836 63384
rect 239680 63096 239732 63102
rect 239680 63038 239732 63044
rect 238760 62824 238812 62830
rect 238760 62766 238812 62772
rect 240796 3534 240824 63378
rect 241428 63096 241480 63102
rect 241428 63038 241480 63044
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 238116 3324 238168 3330
rect 238116 3266 238168 3272
rect 238668 3324 238720 3330
rect 238668 3266 238720 3272
rect 238128 480 238156 3266
rect 239324 480 239352 3470
rect 241440 3466 241468 63038
rect 241624 62966 241652 65484
rect 242636 63238 242664 65484
rect 243556 63374 243584 65484
rect 243544 63368 243596 63374
rect 243544 63310 243596 63316
rect 244188 63368 244240 63374
rect 244188 63310 244240 63316
rect 242624 63232 242676 63238
rect 242624 63174 242676 63180
rect 241612 62960 241664 62966
rect 241612 62902 241664 62908
rect 242808 62960 242860 62966
rect 242808 62902 242860 62908
rect 242820 3534 242848 62902
rect 244096 62824 244148 62830
rect 244096 62766 244148 62772
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 240508 3460 240560 3466
rect 240508 3402 240560 3408
rect 241428 3460 241480 3466
rect 241428 3402 241480 3408
rect 240520 480 240548 3402
rect 241716 480 241744 3470
rect 242912 480 242940 3470
rect 244108 480 244136 62766
rect 244200 3534 244228 63310
rect 244568 62898 244596 65484
rect 244556 62892 244608 62898
rect 244556 62834 244608 62840
rect 245488 62762 245516 65484
rect 246500 63306 246528 65484
rect 246488 63300 246540 63306
rect 246488 63242 246540 63248
rect 246948 63232 247000 63238
rect 246948 63174 247000 63180
rect 245568 62892 245620 62898
rect 245568 62834 245620 62840
rect 245476 62756 245528 62762
rect 245476 62698 245528 62704
rect 245580 6914 245608 62834
rect 245212 6886 245608 6914
rect 244188 3528 244240 3534
rect 244188 3470 244240 3476
rect 245212 480 245240 6886
rect 246960 3534 246988 63174
rect 247420 63170 247448 65484
rect 248328 63504 248380 63510
rect 248328 63446 248380 63452
rect 247408 63164 247460 63170
rect 247408 63106 247460 63112
rect 248340 3534 248368 63446
rect 248432 63034 248460 65484
rect 249352 63442 249380 65484
rect 249340 63436 249392 63442
rect 249340 63378 249392 63384
rect 250364 63102 250392 65484
rect 250352 63096 250404 63102
rect 250352 63038 250404 63044
rect 251088 63096 251140 63102
rect 251088 63038 251140 63044
rect 248420 63028 248472 63034
rect 248420 62970 248472 62976
rect 249708 62280 249760 62286
rect 249708 62222 249760 62228
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 248328 3528 248380 3534
rect 248328 3470 248380 3476
rect 246408 480 246436 3470
rect 247604 480 247632 3470
rect 249720 3466 249748 62222
rect 251100 3534 251128 63038
rect 251284 62966 251312 65484
rect 252296 63374 252324 65484
rect 252284 63368 252336 63374
rect 252284 63310 252336 63316
rect 251272 62960 251324 62966
rect 251272 62902 251324 62908
rect 253216 62830 253244 65484
rect 254228 62898 254256 65484
rect 255148 63238 255176 65484
rect 256160 63510 256188 65484
rect 256148 63504 256200 63510
rect 256148 63446 256200 63452
rect 255136 63232 255188 63238
rect 255136 63174 255188 63180
rect 255964 63164 256016 63170
rect 255964 63106 256016 63112
rect 254216 62892 254268 62898
rect 254216 62834 254268 62840
rect 253204 62824 253256 62830
rect 253204 62766 253256 62772
rect 253848 62824 253900 62830
rect 253848 62766 253900 62772
rect 252376 62212 252428 62218
rect 252376 62154 252428 62160
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 248788 3460 248840 3466
rect 248788 3402 248840 3408
rect 249708 3460 249760 3466
rect 249708 3402 249760 3408
rect 248800 480 248828 3402
rect 249996 480 250024 3470
rect 251192 480 251220 3470
rect 252388 480 252416 62154
rect 252468 62144 252520 62150
rect 252468 62086 252520 62092
rect 252480 3534 252508 62086
rect 253860 6914 253888 62766
rect 253492 6886 253888 6914
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 253492 480 253520 6886
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 254676 3460 254728 3466
rect 254676 3402 254728 3408
rect 254688 480 254716 3402
rect 255884 480 255912 3470
rect 255976 3466 256004 63106
rect 256608 62892 256660 62898
rect 256608 62834 256660 62840
rect 256620 3534 256648 62834
rect 257080 62286 257108 65484
rect 258092 63102 258120 65484
rect 258080 63096 258132 63102
rect 258080 63038 258132 63044
rect 257988 63028 258040 63034
rect 257988 62970 258040 62976
rect 257068 62280 257120 62286
rect 257068 62222 257120 62228
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 255964 3460 256016 3466
rect 255964 3402 256016 3408
rect 258000 3330 258028 62970
rect 259012 62150 259040 65484
rect 259368 62348 259420 62354
rect 259368 62290 259420 62296
rect 259000 62144 259052 62150
rect 259000 62086 259052 62092
rect 259380 3534 259408 62290
rect 260024 62218 260052 65484
rect 260944 62830 260972 65484
rect 261956 63170 261984 65484
rect 261944 63164 261996 63170
rect 261944 63106 261996 63112
rect 262876 62898 262904 65484
rect 263888 63034 263916 65484
rect 263876 63028 263928 63034
rect 263876 62970 263928 62976
rect 262864 62892 262916 62898
rect 262864 62834 262916 62840
rect 260932 62824 260984 62830
rect 260932 62766 260984 62772
rect 260748 62416 260800 62422
rect 260748 62358 260800 62364
rect 260012 62212 260064 62218
rect 260012 62154 260064 62160
rect 260656 62144 260708 62150
rect 260656 62086 260708 62092
rect 260668 16574 260696 62086
rect 260576 16546 260696 16574
rect 260576 3534 260604 16546
rect 260760 6914 260788 62358
rect 264808 62354 264836 65484
rect 264796 62348 264848 62354
rect 264796 62290 264848 62296
rect 263508 62280 263560 62286
rect 263508 62222 263560 62228
rect 260668 6886 260788 6914
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 260564 3528 260616 3534
rect 260564 3470 260616 3476
rect 257068 3324 257120 3330
rect 257068 3266 257120 3272
rect 257988 3324 258040 3330
rect 257988 3266 258040 3272
rect 257080 480 257108 3266
rect 258276 480 258304 3470
rect 259472 480 259500 3470
rect 260668 480 260696 6886
rect 263520 3534 263548 62222
rect 264888 62212 264940 62218
rect 264888 62154 264940 62160
rect 264900 3534 264928 62154
rect 265820 62150 265848 65484
rect 266740 62422 266768 65484
rect 267648 63096 267700 63102
rect 267648 63038 267700 63044
rect 267004 62960 267056 62966
rect 267004 62902 267056 62908
rect 266728 62416 266780 62422
rect 266728 62358 266780 62364
rect 265808 62144 265860 62150
rect 265808 62086 265860 62092
rect 267016 3534 267044 62902
rect 267096 62144 267148 62150
rect 267096 62086 267148 62092
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 267004 3528 267056 3534
rect 267004 3470 267056 3476
rect 261760 3324 261812 3330
rect 261760 3266 261812 3272
rect 261772 480 261800 3266
rect 262968 480 262996 3470
rect 264164 480 264192 3470
rect 265360 480 265388 3470
rect 266544 3460 266596 3466
rect 266544 3402 266596 3408
rect 266556 480 266584 3402
rect 267108 3330 267136 62086
rect 267660 3466 267688 63038
rect 267752 62150 267780 65484
rect 268672 62286 268700 65484
rect 269028 62348 269080 62354
rect 269028 62290 269080 62296
rect 268660 62280 268712 62286
rect 268660 62222 268712 62228
rect 267740 62144 267792 62150
rect 267740 62086 267792 62092
rect 269040 6914 269068 62290
rect 269684 62218 269712 65484
rect 270604 62966 270632 65484
rect 271616 63102 271644 65484
rect 271604 63096 271656 63102
rect 271604 63038 271656 63044
rect 270592 62960 270644 62966
rect 270592 62902 270644 62908
rect 270408 62280 270460 62286
rect 270408 62222 270460 62228
rect 269672 62212 269724 62218
rect 269672 62154 269724 62160
rect 269764 62144 269816 62150
rect 269764 62086 269816 62092
rect 268856 6886 269068 6914
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 267096 3324 267148 3330
rect 267096 3266 267148 3272
rect 267752 480 267780 3470
rect 268856 480 268884 6886
rect 269776 3534 269804 62086
rect 270420 6914 270448 62222
rect 271788 62212 271840 62218
rect 271788 62154 271840 62160
rect 270052 6886 270448 6914
rect 269764 3528 269816 3534
rect 269764 3470 269816 3476
rect 270052 480 270080 6886
rect 271800 3534 271828 62154
rect 272536 62150 272564 65484
rect 273548 62354 273576 65484
rect 273536 62348 273588 62354
rect 273536 62290 273588 62296
rect 274468 62286 274496 65484
rect 274456 62280 274508 62286
rect 274456 62222 274508 62228
rect 274548 62280 274600 62286
rect 274548 62222 274600 62228
rect 272524 62144 272576 62150
rect 272524 62086 272576 62092
rect 274560 3534 274588 62222
rect 275480 62218 275508 65484
rect 275468 62212 275520 62218
rect 275468 62154 275520 62160
rect 275928 62212 275980 62218
rect 275928 62154 275980 62160
rect 275940 3534 275968 62154
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 275928 3528 275980 3534
rect 275928 3470 275980 3476
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 271248 480 271276 3470
rect 272432 3324 272484 3330
rect 272432 3266 272484 3272
rect 272444 480 272472 3266
rect 273640 480 273668 3470
rect 274836 480 274864 3470
rect 276032 480 276060 3470
rect 276400 3330 276428 65484
rect 277216 62824 277268 62830
rect 277216 62766 277268 62772
rect 277228 6914 277256 62766
rect 277412 62286 277440 65484
rect 277400 62280 277452 62286
rect 277400 62222 277452 62228
rect 278332 62218 278360 65484
rect 278320 62212 278372 62218
rect 278320 62154 278372 62160
rect 278688 62212 278740 62218
rect 278688 62154 278740 62160
rect 277308 62144 277360 62150
rect 277308 62086 277360 62092
rect 277136 6886 277256 6914
rect 276388 3324 276440 3330
rect 276388 3266 276440 3272
rect 277136 480 277164 6886
rect 277320 3534 277348 62086
rect 278700 6914 278728 62154
rect 279344 62150 279372 65484
rect 280264 62830 280292 65484
rect 280252 62824 280304 62830
rect 280252 62766 280304 62772
rect 281276 62218 281304 65484
rect 281264 62212 281316 62218
rect 281264 62154 281316 62160
rect 281448 62212 281500 62218
rect 281448 62154 281500 62160
rect 279332 62144 279384 62150
rect 279332 62086 279384 62092
rect 280804 62144 280856 62150
rect 280804 62086 280856 62092
rect 278332 6886 278728 6914
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 278332 480 278360 6886
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 279516 3324 279568 3330
rect 279516 3266 279568 3272
rect 279528 480 279556 3266
rect 280724 480 280752 3470
rect 280816 3330 280844 62086
rect 281460 3534 281488 62154
rect 282196 62150 282224 65484
rect 283208 62218 283236 65484
rect 283196 62212 283248 62218
rect 283196 62154 283248 62160
rect 284128 62150 284156 65484
rect 282184 62144 282236 62150
rect 282184 62086 282236 62092
rect 282828 62144 282880 62150
rect 282828 62086 282880 62092
rect 284116 62144 284168 62150
rect 284116 62086 284168 62092
rect 282840 3534 282868 62086
rect 285140 3534 285168 65484
rect 285588 62144 285640 62150
rect 285588 62086 285640 62092
rect 285600 6914 285628 62086
rect 285416 6886 285628 6914
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281908 3528 281960 3534
rect 281908 3470 281960 3476
rect 282828 3528 282880 3534
rect 282828 3470 282880 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 285128 3528 285180 3534
rect 285128 3470 285180 3476
rect 280804 3324 280856 3330
rect 280804 3266 280856 3272
rect 281920 480 281948 3470
rect 283116 480 283144 3470
rect 284300 2984 284352 2990
rect 284300 2926 284352 2932
rect 284312 480 284340 2926
rect 285416 480 285444 6886
rect 286060 2990 286088 65484
rect 287072 62150 287100 65484
rect 287060 62144 287112 62150
rect 287060 62086 287112 62092
rect 287992 3466 288020 65484
rect 289004 62150 289032 65484
rect 289924 64874 289952 65484
rect 289832 64846 289952 64874
rect 289832 62234 289860 64846
rect 289740 62206 289860 62234
rect 288348 62144 288400 62150
rect 288348 62086 288400 62092
rect 288992 62144 289044 62150
rect 288992 62086 289044 62092
rect 286600 3460 286652 3466
rect 286600 3402 286652 3408
rect 287980 3460 288032 3466
rect 287980 3402 288032 3408
rect 286048 2984 286100 2990
rect 286048 2926 286100 2932
rect 286612 480 286640 3402
rect 288360 2922 288388 62086
rect 289740 3534 289768 62206
rect 290936 62150 290964 65484
rect 289820 62144 289872 62150
rect 289820 62086 289872 62092
rect 290924 62144 290976 62150
rect 290924 62086 290976 62092
rect 289832 16574 289860 62086
rect 289832 16546 290228 16574
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 287796 2916 287848 2922
rect 287796 2858 287848 2864
rect 288348 2916 288400 2922
rect 288348 2858 288400 2864
rect 287808 480 287836 2858
rect 289004 480 289032 3470
rect 290200 480 290228 16546
rect 291856 3534 291884 65484
rect 292580 62144 292632 62150
rect 292580 62086 292632 62092
rect 292592 11762 292620 62086
rect 292580 11756 292632 11762
rect 292580 11698 292632 11704
rect 292868 6914 292896 65484
rect 293788 62150 293816 65484
rect 293776 62144 293828 62150
rect 293776 62086 293828 62092
rect 294800 16574 294828 65484
rect 295720 16574 295748 65484
rect 296732 16574 296760 65484
rect 297652 62150 297680 65484
rect 298664 62150 298692 65484
rect 299584 64874 299612 65484
rect 300596 64874 300624 65484
rect 299584 64846 299704 64874
rect 300596 64846 300808 64874
rect 297640 62144 297692 62150
rect 297640 62086 297692 62092
rect 298192 62144 298244 62150
rect 298192 62086 298244 62092
rect 298652 62144 298704 62150
rect 298652 62086 298704 62092
rect 299388 62144 299440 62150
rect 299388 62086 299440 62092
rect 298204 16574 298232 62086
rect 294800 16546 294920 16574
rect 295720 16546 296116 16574
rect 296732 16546 297312 16574
rect 298204 16546 298508 16574
rect 293684 11756 293736 11762
rect 293684 11698 293736 11704
rect 292592 6886 292896 6914
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291844 3528 291896 3534
rect 291844 3470 291896 3476
rect 291396 480 291424 3470
rect 292592 480 292620 6886
rect 293696 480 293724 11698
rect 294892 480 294920 16546
rect 296088 480 296116 16546
rect 297284 480 297312 16546
rect 298480 480 298508 16546
rect 299400 3482 299428 62086
rect 299676 16574 299704 64846
rect 299676 16546 300716 16574
rect 300688 3482 300716 16546
rect 300780 3602 300808 64846
rect 301516 62150 301544 65484
rect 302528 62762 302556 65484
rect 303448 64874 303476 65484
rect 303448 64846 303568 64874
rect 302516 62756 302568 62762
rect 302516 62698 302568 62704
rect 303344 62756 303396 62762
rect 303344 62698 303396 62704
rect 301504 62144 301556 62150
rect 301504 62086 301556 62092
rect 302424 62144 302476 62150
rect 302424 62086 302476 62092
rect 302436 16574 302464 62086
rect 302436 16546 303200 16574
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 301964 3596 302016 3602
rect 301964 3538 302016 3544
rect 299400 3454 299704 3482
rect 300688 3454 300808 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3454
rect 301976 480 302004 3538
rect 303172 480 303200 16546
rect 303356 3534 303384 62698
rect 303540 3602 303568 64846
rect 304460 62150 304488 65484
rect 305380 62150 305408 65484
rect 306392 62150 306420 65484
rect 307312 64874 307340 65484
rect 307312 64846 307616 64874
rect 304448 62144 304500 62150
rect 304448 62086 304500 62092
rect 304908 62144 304960 62150
rect 304908 62086 304960 62092
rect 305368 62144 305420 62150
rect 305368 62086 305420 62092
rect 306288 62144 306340 62150
rect 306288 62086 306340 62092
rect 306380 62144 306432 62150
rect 306380 62086 306432 62092
rect 303528 3596 303580 3602
rect 303528 3538 303580 3544
rect 303344 3528 303396 3534
rect 303344 3470 303396 3476
rect 304356 3528 304408 3534
rect 304356 3470 304408 3476
rect 304368 480 304396 3470
rect 304920 3466 304948 62086
rect 305552 3596 305604 3602
rect 305552 3538 305604 3544
rect 304908 3460 304960 3466
rect 304908 3402 304960 3408
rect 305564 480 305592 3538
rect 306300 3330 306328 62086
rect 307588 3466 307616 64846
rect 308324 62422 308352 65484
rect 308312 62416 308364 62422
rect 308312 62358 308364 62364
rect 309244 62150 309272 65484
rect 310256 64874 310284 65484
rect 310256 64846 310468 64874
rect 309784 62416 309836 62422
rect 309784 62358 309836 62364
rect 307668 62144 307720 62150
rect 307668 62086 307720 62092
rect 309232 62144 309284 62150
rect 309232 62086 309284 62092
rect 307680 3534 307708 62086
rect 309796 3534 309824 62358
rect 310336 62144 310388 62150
rect 310336 62086 310388 62092
rect 307668 3528 307720 3534
rect 307668 3470 307720 3476
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 306748 3460 306800 3466
rect 306748 3402 306800 3408
rect 307576 3460 307628 3466
rect 307576 3402 307628 3408
rect 306288 3324 306340 3330
rect 306288 3266 306340 3272
rect 306760 480 306788 3402
rect 307944 3324 307996 3330
rect 307944 3266 307996 3272
rect 307956 480 307984 3266
rect 309060 480 309088 3470
rect 310244 3460 310296 3466
rect 310244 3402 310296 3408
rect 310256 480 310284 3402
rect 310348 3194 310376 62086
rect 310440 3602 310468 64846
rect 311176 63034 311204 65484
rect 311164 63028 311216 63034
rect 311164 62970 311216 62976
rect 311808 63028 311860 63034
rect 311808 62970 311860 62976
rect 310428 3596 310480 3602
rect 310428 3538 310480 3544
rect 311820 3534 311848 62970
rect 312188 62150 312216 65484
rect 313108 62694 313136 65484
rect 313096 62688 313148 62694
rect 313096 62630 313148 62636
rect 313924 62688 313976 62694
rect 313924 62630 313976 62636
rect 312176 62144 312228 62150
rect 312176 62086 312228 62092
rect 313188 62144 313240 62150
rect 313188 62086 313240 62092
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 311808 3528 311860 3534
rect 311808 3470 311860 3476
rect 310336 3188 310388 3194
rect 310336 3130 310388 3136
rect 311452 480 311480 3470
rect 312636 3188 312688 3194
rect 312636 3130 312688 3136
rect 312648 480 312676 3130
rect 313200 3126 313228 62086
rect 313832 3596 313884 3602
rect 313832 3538 313884 3544
rect 313188 3120 313240 3126
rect 313188 3062 313240 3068
rect 313844 480 313872 3538
rect 313936 3398 313964 62630
rect 314120 62150 314148 65484
rect 315040 62218 315068 65484
rect 316052 62354 316080 65484
rect 316972 64874 317000 65484
rect 316972 64846 317276 64874
rect 316040 62348 316092 62354
rect 316040 62290 316092 62296
rect 315028 62212 315080 62218
rect 315028 62154 315080 62160
rect 314108 62144 314160 62150
rect 314108 62086 314160 62092
rect 314568 62144 314620 62150
rect 314568 62086 314620 62092
rect 314580 3874 314608 62086
rect 314568 3868 314620 3874
rect 314568 3810 314620 3816
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 313924 3392 313976 3398
rect 313924 3334 313976 3340
rect 315040 480 315068 3470
rect 317248 3194 317276 64846
rect 317328 62348 317380 62354
rect 317328 62290 317380 62296
rect 317340 3602 317368 62290
rect 317984 62150 318012 65484
rect 318904 63034 318932 65484
rect 318892 63028 318944 63034
rect 318892 62970 318944 62976
rect 319916 62286 319944 65484
rect 319904 62280 319956 62286
rect 319904 62222 319956 62228
rect 318064 62212 318116 62218
rect 318064 62154 318116 62160
rect 317972 62144 318024 62150
rect 317972 62086 318024 62092
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 318076 3534 318104 62154
rect 320836 62150 320864 65484
rect 321008 63028 321060 63034
rect 321008 62970 321060 62976
rect 320916 62280 320968 62286
rect 320916 62222 320968 62228
rect 318708 62144 318760 62150
rect 318708 62086 318760 62092
rect 320824 62144 320876 62150
rect 320824 62086 320876 62092
rect 318524 3868 318576 3874
rect 318524 3810 318576 3816
rect 318064 3528 318116 3534
rect 318064 3470 318116 3476
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317236 3188 317288 3194
rect 317236 3130 317288 3136
rect 316224 3120 316276 3126
rect 316224 3062 316276 3068
rect 316236 480 316264 3062
rect 317340 480 317368 3334
rect 318536 480 318564 3810
rect 318720 3262 318748 62086
rect 320928 3738 320956 62222
rect 320916 3732 320968 3738
rect 320916 3674 320968 3680
rect 320916 3596 320968 3602
rect 320916 3538 320968 3544
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 318708 3256 318760 3262
rect 318708 3198 318760 3204
rect 319732 480 319760 3470
rect 320928 480 320956 3538
rect 321020 3330 321048 62970
rect 321848 62490 321876 65484
rect 321836 62484 321888 62490
rect 321836 62426 321888 62432
rect 321468 62144 321520 62150
rect 321468 62086 321520 62092
rect 321008 3324 321060 3330
rect 321008 3266 321060 3272
rect 321480 3058 321508 62086
rect 322768 3466 322796 65484
rect 322848 62484 322900 62490
rect 322848 62426 322900 62432
rect 322860 4146 322888 62426
rect 323780 62150 323808 65484
rect 324700 62150 324728 65484
rect 325712 62762 325740 65484
rect 326632 64874 326660 65484
rect 326632 64846 327028 64874
rect 325700 62756 325752 62762
rect 325700 62698 325752 62704
rect 323768 62144 323820 62150
rect 323768 62086 323820 62092
rect 324228 62144 324280 62150
rect 324228 62086 324280 62092
rect 324688 62144 324740 62150
rect 324688 62086 324740 62092
rect 325608 62144 325660 62150
rect 325608 62086 325660 62092
rect 322848 4140 322900 4146
rect 322848 4082 322900 4088
rect 324240 3670 324268 62086
rect 325620 3738 325648 62086
rect 325516 3732 325568 3738
rect 325516 3674 325568 3680
rect 325608 3732 325660 3738
rect 325608 3674 325660 3680
rect 324228 3664 324280 3670
rect 324228 3606 324280 3612
rect 325528 3482 325556 3674
rect 322756 3460 322808 3466
rect 325528 3454 325648 3482
rect 322756 3402 322808 3408
rect 324412 3324 324464 3330
rect 324412 3266 324464 3272
rect 323308 3256 323360 3262
rect 323308 3198 323360 3204
rect 322112 3188 322164 3194
rect 322112 3130 322164 3136
rect 321468 3052 321520 3058
rect 321468 2994 321520 3000
rect 322124 480 322152 3130
rect 323320 480 323348 3198
rect 324424 480 324452 3266
rect 325620 480 325648 3454
rect 326804 3052 326856 3058
rect 326804 2994 326856 3000
rect 326816 480 326844 2994
rect 327000 2990 327028 64846
rect 327644 62898 327672 65484
rect 328564 63170 328592 65484
rect 329576 64874 329604 65484
rect 329576 64846 329788 64874
rect 328552 63164 328604 63170
rect 328552 63106 328604 63112
rect 329656 63164 329708 63170
rect 329656 63106 329708 63112
rect 327632 62892 327684 62898
rect 327632 62834 327684 62840
rect 328368 62892 328420 62898
rect 328368 62834 328420 62840
rect 328000 4140 328052 4146
rect 328000 4082 328052 4088
rect 326988 2984 327040 2990
rect 326988 2926 327040 2932
rect 328012 480 328040 4082
rect 328380 3330 328408 62834
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 328368 3324 328420 3330
rect 328368 3266 328420 3272
rect 329208 480 329236 3402
rect 329668 3194 329696 63106
rect 329656 3188 329708 3194
rect 329656 3130 329708 3136
rect 329760 3058 329788 64846
rect 330496 63034 330524 65484
rect 330484 63028 330536 63034
rect 330484 62970 330536 62976
rect 331128 63028 331180 63034
rect 331128 62970 331180 62976
rect 331140 3670 331168 62970
rect 331508 62150 331536 65484
rect 332428 64874 332456 65484
rect 332428 64846 332548 64874
rect 331864 62756 331916 62762
rect 331864 62698 331916 62704
rect 331496 62144 331548 62150
rect 331496 62086 331548 62092
rect 331588 3732 331640 3738
rect 331588 3674 331640 3680
rect 330392 3664 330444 3670
rect 330392 3606 330444 3612
rect 331128 3664 331180 3670
rect 331128 3606 331180 3612
rect 329748 3052 329800 3058
rect 329748 2994 329800 3000
rect 330404 480 330432 3606
rect 331600 480 331628 3674
rect 331876 3534 331904 62698
rect 332324 62144 332376 62150
rect 332324 62086 332376 62092
rect 332336 3738 332364 62086
rect 332324 3732 332376 3738
rect 332324 3674 332376 3680
rect 331864 3528 331916 3534
rect 331864 3470 331916 3476
rect 332520 3466 332548 64846
rect 333440 62490 333468 65484
rect 334360 63374 334388 65484
rect 334348 63368 334400 63374
rect 334348 63310 334400 63316
rect 335268 63368 335320 63374
rect 335268 63310 335320 63316
rect 333428 62484 333480 62490
rect 333428 62426 333480 62432
rect 334624 62484 334676 62490
rect 334624 62426 334676 62432
rect 334636 4010 334664 62426
rect 334624 4004 334676 4010
rect 334624 3946 334676 3952
rect 335280 3806 335308 63310
rect 335372 62354 335400 65484
rect 336292 64874 336320 65484
rect 336292 64846 336596 64874
rect 335360 62348 335412 62354
rect 335360 62290 335412 62296
rect 336568 3874 336596 64846
rect 336648 62348 336700 62354
rect 336648 62290 336700 62296
rect 336556 3868 336608 3874
rect 336556 3810 336608 3816
rect 335268 3800 335320 3806
rect 335268 3742 335320 3748
rect 336660 3602 336688 62290
rect 337304 62150 337332 65484
rect 338224 62354 338252 65484
rect 339236 64874 339264 65484
rect 339236 64846 339356 64874
rect 338212 62348 338264 62354
rect 338212 62290 338264 62296
rect 337292 62144 337344 62150
rect 337292 62086 337344 62092
rect 338672 3664 338724 3670
rect 338672 3606 338724 3612
rect 336648 3596 336700 3602
rect 336648 3538 336700 3544
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 332508 3460 332560 3466
rect 332508 3402 332560 3408
rect 332704 480 332732 3470
rect 335084 3324 335136 3330
rect 335084 3266 335136 3272
rect 333888 2984 333940 2990
rect 333888 2926 333940 2932
rect 333900 480 333928 2926
rect 335096 480 335124 3266
rect 336280 3188 336332 3194
rect 336280 3130 336332 3136
rect 336292 480 336320 3130
rect 337476 3052 337528 3058
rect 337476 2994 337528 3000
rect 337488 480 337516 2994
rect 338684 480 338712 3606
rect 339328 3534 339356 64846
rect 340156 62830 340184 65484
rect 340144 62824 340196 62830
rect 340144 62766 340196 62772
rect 340788 62824 340840 62830
rect 340788 62766 340840 62772
rect 339408 62348 339460 62354
rect 339408 62290 339460 62296
rect 339420 3670 339448 62290
rect 340236 62144 340288 62150
rect 340236 62086 340288 62092
rect 339868 3732 339920 3738
rect 339868 3674 339920 3680
rect 339408 3664 339460 3670
rect 339408 3606 339460 3612
rect 339316 3528 339368 3534
rect 339316 3470 339368 3476
rect 339880 480 339908 3674
rect 340248 3126 340276 62086
rect 340800 3738 340828 62766
rect 341168 62422 341196 65484
rect 341156 62416 341208 62422
rect 341156 62358 341208 62364
rect 340788 3732 340840 3738
rect 340788 3674 340840 3680
rect 342088 3466 342116 65484
rect 342168 62416 342220 62422
rect 342168 62358 342220 62364
rect 342180 4146 342208 62358
rect 343100 62150 343128 65484
rect 344020 62150 344048 65484
rect 345032 62150 345060 65484
rect 345952 64874 345980 65484
rect 345952 64846 346348 64874
rect 343088 62144 343140 62150
rect 343088 62086 343140 62092
rect 343548 62144 343600 62150
rect 343548 62086 343600 62092
rect 344008 62144 344060 62150
rect 344008 62086 344060 62092
rect 344928 62144 344980 62150
rect 344928 62086 344980 62092
rect 345020 62144 345072 62150
rect 345020 62086 345072 62092
rect 346216 62144 346268 62150
rect 346216 62086 346268 62092
rect 342168 4140 342220 4146
rect 342168 4082 342220 4088
rect 343560 4010 343588 62086
rect 344940 4078 344968 62086
rect 344928 4072 344980 4078
rect 344928 4014 344980 4020
rect 342168 4004 342220 4010
rect 342168 3946 342220 3952
rect 343548 4004 343600 4010
rect 343548 3946 343600 3952
rect 340972 3460 341024 3466
rect 340972 3402 341024 3408
rect 342076 3460 342128 3466
rect 342076 3402 342128 3408
rect 340236 3120 340288 3126
rect 340236 3062 340288 3068
rect 340984 480 341012 3402
rect 342180 480 342208 3946
rect 346228 3874 346256 62086
rect 346216 3868 346268 3874
rect 346216 3810 346268 3816
rect 343364 3800 343416 3806
rect 343364 3742 343416 3748
rect 343376 480 343404 3742
rect 346320 3602 346348 64846
rect 346964 62898 346992 65484
rect 346952 62892 347004 62898
rect 346952 62834 347004 62840
rect 347688 62892 347740 62898
rect 347688 62834 347740 62840
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 345756 3596 345808 3602
rect 345756 3538 345808 3544
rect 346308 3596 346360 3602
rect 346308 3538 346360 3544
rect 344572 480 344600 3538
rect 345768 480 345796 3538
rect 347700 3330 347728 62834
rect 347884 62150 347912 65484
rect 348896 64874 348924 65484
rect 348896 64846 349016 64874
rect 347872 62144 347924 62150
rect 347872 62086 347924 62092
rect 348988 3670 349016 64846
rect 349816 63034 349844 65484
rect 349804 63028 349856 63034
rect 349804 62970 349856 62976
rect 350448 63028 350500 63034
rect 350448 62970 350500 62976
rect 349068 62144 349120 62150
rect 349068 62086 349120 62092
rect 349080 3942 349108 62086
rect 350460 6914 350488 62970
rect 350828 62150 350856 65484
rect 351748 62694 351776 65484
rect 351736 62688 351788 62694
rect 351736 62630 351788 62636
rect 352564 62688 352616 62694
rect 352564 62630 352616 62636
rect 350816 62144 350868 62150
rect 350816 62086 350868 62092
rect 351828 62144 351880 62150
rect 351828 62086 351880 62092
rect 350368 6886 350488 6914
rect 349068 3936 349120 3942
rect 349068 3878 349120 3884
rect 350368 3806 350396 6886
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 350356 3800 350408 3806
rect 350356 3742 350408 3748
rect 350448 3732 350500 3738
rect 350448 3674 350500 3680
rect 348056 3664 348108 3670
rect 348056 3606 348108 3612
rect 348976 3664 349028 3670
rect 348976 3606 349028 3612
rect 347688 3324 347740 3330
rect 347688 3266 347740 3272
rect 346952 3120 347004 3126
rect 346952 3062 347004 3068
rect 346964 480 346992 3062
rect 348068 480 348096 3606
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 349264 480 349292 3470
rect 350460 480 350488 3674
rect 351656 480 351684 4082
rect 351840 3398 351868 62086
rect 352576 3534 352604 62630
rect 352760 62150 352788 65484
rect 353680 63374 353708 65484
rect 353668 63368 353720 63374
rect 353668 63310 353720 63316
rect 354588 63368 354640 63374
rect 354588 63310 354640 63316
rect 352748 62144 352800 62150
rect 352748 62086 352800 62092
rect 353208 62144 353260 62150
rect 353208 62086 353260 62092
rect 353220 3738 353248 62086
rect 354036 4004 354088 4010
rect 354036 3946 354088 3952
rect 353208 3732 353260 3738
rect 353208 3674 353260 3680
rect 352564 3528 352616 3534
rect 352564 3470 352616 3476
rect 352840 3460 352892 3466
rect 352840 3402 352892 3408
rect 351828 3392 351880 3398
rect 351828 3334 351880 3340
rect 352852 480 352880 3402
rect 354048 480 354076 3946
rect 354600 3262 354628 63310
rect 354692 62150 354720 65484
rect 355612 64874 355640 65484
rect 355612 64846 356008 64874
rect 354680 62144 354732 62150
rect 354680 62086 354732 62092
rect 355876 62144 355928 62150
rect 355876 62086 355928 62092
rect 355888 4146 355916 62086
rect 355876 4140 355928 4146
rect 355876 4082 355928 4088
rect 355232 4072 355284 4078
rect 355232 4014 355284 4020
rect 354588 3256 354640 3262
rect 354588 3198 354640 3204
rect 355244 480 355272 4014
rect 355980 4010 356008 64846
rect 356624 62150 356652 65484
rect 357544 62354 357572 65484
rect 358556 64874 358584 65484
rect 358556 64846 358676 64874
rect 357532 62348 357584 62354
rect 357532 62290 357584 62296
rect 356612 62144 356664 62150
rect 356612 62086 356664 62092
rect 357348 62144 357400 62150
rect 357348 62086 357400 62092
rect 355968 4004 356020 4010
rect 355968 3946 356020 3952
rect 356336 3868 356388 3874
rect 356336 3810 356388 3816
rect 356348 480 356376 3810
rect 357360 3466 357388 62086
rect 358648 3602 358676 64846
rect 359476 62830 359504 65484
rect 359464 62824 359516 62830
rect 359464 62766 359516 62772
rect 360108 62824 360160 62830
rect 360108 62766 360160 62772
rect 358728 62348 358780 62354
rect 358728 62290 358780 62296
rect 358740 4078 358768 62290
rect 358728 4072 358780 4078
rect 358728 4014 358780 4020
rect 359924 3936 359976 3942
rect 359924 3878 359976 3884
rect 357532 3596 357584 3602
rect 357532 3538 357584 3544
rect 358636 3596 358688 3602
rect 358636 3538 358688 3544
rect 357348 3460 357400 3466
rect 357348 3402 357400 3408
rect 357544 480 357572 3538
rect 358728 3324 358780 3330
rect 358728 3266 358780 3272
rect 358740 480 358768 3266
rect 359936 480 359964 3878
rect 360120 3874 360148 62766
rect 360488 62422 360516 65484
rect 360476 62416 360528 62422
rect 360476 62358 360528 62364
rect 360108 3868 360160 3874
rect 360108 3810 360160 3816
rect 361408 3670 361436 65484
rect 361488 62416 361540 62422
rect 361488 62358 361540 62364
rect 361120 3664 361172 3670
rect 361120 3606 361172 3612
rect 361396 3664 361448 3670
rect 361396 3606 361448 3612
rect 361132 480 361160 3606
rect 361500 3330 361528 62358
rect 362420 62150 362448 65484
rect 363340 62150 363368 65484
rect 364352 62150 364380 65484
rect 365272 64874 365300 65484
rect 365272 64846 365576 64874
rect 362408 62144 362460 62150
rect 362408 62086 362460 62092
rect 362868 62144 362920 62150
rect 362868 62086 362920 62092
rect 363328 62144 363380 62150
rect 363328 62086 363380 62092
rect 364248 62144 364300 62150
rect 364248 62086 364300 62092
rect 364340 62144 364392 62150
rect 364340 62086 364392 62092
rect 362880 3942 362908 62086
rect 362868 3936 362920 3942
rect 362868 3878 362920 3884
rect 362316 3800 362368 3806
rect 362316 3742 362368 3748
rect 361488 3324 361540 3330
rect 361488 3266 361540 3272
rect 362328 480 362356 3742
rect 363512 3392 363564 3398
rect 363512 3334 363564 3340
rect 363524 480 363552 3334
rect 364260 2922 364288 62086
rect 365548 3534 365576 64846
rect 366284 62898 366312 65484
rect 367204 63170 367232 65484
rect 368216 64874 368244 65484
rect 368216 64846 368428 64874
rect 367192 63164 367244 63170
rect 367192 63106 367244 63112
rect 368296 63164 368348 63170
rect 368296 63106 368348 63112
rect 366272 62892 366324 62898
rect 366272 62834 366324 62840
rect 367008 62892 367060 62898
rect 367008 62834 367060 62840
rect 365628 62144 365680 62150
rect 365628 62086 365680 62092
rect 364616 3528 364668 3534
rect 364616 3470 364668 3476
rect 365536 3528 365588 3534
rect 365536 3470 365588 3476
rect 364248 2916 364300 2922
rect 364248 2858 364300 2864
rect 364628 480 364656 3470
rect 365640 2990 365668 62086
rect 367020 3806 367048 62834
rect 368204 4140 368256 4146
rect 368204 4082 368256 4088
rect 367008 3800 367060 3806
rect 367008 3742 367060 3748
rect 365812 3732 365864 3738
rect 365812 3674 365864 3680
rect 365628 2984 365680 2990
rect 365628 2926 365680 2932
rect 365824 480 365852 3674
rect 367008 3256 367060 3262
rect 367008 3198 367060 3204
rect 367020 480 367048 3198
rect 368216 480 368244 4082
rect 368308 3058 368336 63106
rect 368400 3738 368428 64846
rect 369136 63034 369164 65484
rect 369124 63028 369176 63034
rect 369124 62970 369176 62976
rect 369768 63028 369820 63034
rect 369768 62970 369820 62976
rect 369400 4004 369452 4010
rect 369400 3946 369452 3952
rect 368388 3732 368440 3738
rect 368388 3674 368440 3680
rect 368296 3052 368348 3058
rect 368296 2994 368348 3000
rect 369412 480 369440 3946
rect 369780 3398 369808 62970
rect 370148 62150 370176 65484
rect 370136 62144 370188 62150
rect 370136 62086 370188 62092
rect 371068 3466 371096 65484
rect 372080 62150 372108 65484
rect 373000 63374 373028 65484
rect 372988 63368 373040 63374
rect 372988 63310 373040 63316
rect 373908 63368 373960 63374
rect 373908 63310 373960 63316
rect 371148 62144 371200 62150
rect 371148 62086 371200 62092
rect 372068 62144 372120 62150
rect 372068 62086 372120 62092
rect 372528 62144 372580 62150
rect 372528 62086 372580 62092
rect 370596 3460 370648 3466
rect 370596 3402 370648 3408
rect 371056 3460 371108 3466
rect 371056 3402 371108 3408
rect 369768 3392 369820 3398
rect 369768 3334 369820 3340
rect 370608 480 370636 3402
rect 371160 3126 371188 62086
rect 371700 4072 371752 4078
rect 371700 4014 371752 4020
rect 371148 3120 371200 3126
rect 371148 3062 371200 3068
rect 371712 480 371740 4014
rect 372540 4010 372568 62086
rect 373920 4146 373948 63310
rect 374012 62354 374040 65484
rect 374932 64874 374960 65484
rect 374932 64846 375236 64874
rect 374000 62348 374052 62354
rect 374000 62290 374052 62296
rect 373908 4140 373960 4146
rect 373908 4082 373960 4088
rect 375208 4078 375236 64846
rect 375288 62348 375340 62354
rect 375288 62290 375340 62296
rect 375196 4072 375248 4078
rect 375196 4014 375248 4020
rect 372528 4004 372580 4010
rect 372528 3946 372580 3952
rect 375300 3890 375328 62290
rect 375944 62150 375972 65484
rect 376864 62354 376892 65484
rect 377876 64874 377904 65484
rect 377876 64846 377996 64874
rect 376852 62348 376904 62354
rect 376852 62290 376904 62296
rect 375932 62144 375984 62150
rect 375932 62086 375984 62092
rect 376668 62144 376720 62150
rect 376668 62086 376720 62092
rect 374092 3868 374144 3874
rect 374092 3810 374144 3816
rect 375208 3862 375328 3890
rect 372896 3596 372948 3602
rect 372896 3538 372948 3544
rect 372908 480 372936 3538
rect 374104 480 374132 3810
rect 375208 3262 375236 3862
rect 376484 3664 376536 3670
rect 376484 3606 376536 3612
rect 375288 3324 375340 3330
rect 375288 3266 375340 3272
rect 375196 3256 375248 3262
rect 375196 3198 375248 3204
rect 375300 480 375328 3266
rect 376496 480 376524 3606
rect 376680 3262 376708 62086
rect 377680 3936 377732 3942
rect 377680 3878 377732 3884
rect 376668 3256 376720 3262
rect 376668 3198 376720 3204
rect 377692 480 377720 3878
rect 377968 3602 377996 64846
rect 378796 62830 378824 65484
rect 378784 62824 378836 62830
rect 378784 62766 378836 62772
rect 379428 62824 379480 62830
rect 379428 62766 379480 62772
rect 378048 62348 378100 62354
rect 378048 62290 378100 62296
rect 377956 3596 378008 3602
rect 377956 3538 378008 3544
rect 378060 3194 378088 62290
rect 379440 3942 379468 62766
rect 379808 62354 379836 65484
rect 380728 64874 380756 65484
rect 380728 64846 380848 64874
rect 379796 62348 379848 62354
rect 379796 62290 379848 62296
rect 379428 3936 379480 3942
rect 379428 3878 379480 3884
rect 380820 3874 380848 64846
rect 381544 62348 381596 62354
rect 381544 62290 381596 62296
rect 381556 4826 381584 62290
rect 381740 62150 381768 65484
rect 382660 62150 382688 65484
rect 383672 62150 383700 65484
rect 384592 64874 384620 65484
rect 384592 64846 384988 64874
rect 381728 62144 381780 62150
rect 381728 62086 381780 62092
rect 382188 62144 382240 62150
rect 382188 62086 382240 62092
rect 382648 62144 382700 62150
rect 382648 62086 382700 62092
rect 383568 62144 383620 62150
rect 383568 62086 383620 62092
rect 383660 62144 383712 62150
rect 383660 62086 383712 62092
rect 384856 62144 384908 62150
rect 384856 62086 384908 62092
rect 381544 4820 381596 4826
rect 381544 4762 381596 4768
rect 380808 3868 380860 3874
rect 380808 3810 380860 3816
rect 382200 3670 382228 62086
rect 383580 5234 383608 62086
rect 383568 5228 383620 5234
rect 383568 5170 383620 5176
rect 384868 3806 384896 62086
rect 382372 3800 382424 3806
rect 382372 3742 382424 3748
rect 384856 3800 384908 3806
rect 384856 3742 384908 3748
rect 382188 3664 382240 3670
rect 382188 3606 382240 3612
rect 381176 3528 381228 3534
rect 381176 3470 381228 3476
rect 378048 3188 378100 3194
rect 378048 3130 378100 3136
rect 379980 2984 380032 2990
rect 379980 2926 380032 2932
rect 378876 2916 378928 2922
rect 378876 2858 378928 2864
rect 378888 480 378916 2858
rect 379992 480 380020 2926
rect 381188 480 381216 3470
rect 382384 480 382412 3742
rect 384764 3732 384816 3738
rect 384764 3674 384816 3680
rect 383568 3052 383620 3058
rect 383568 2994 383620 3000
rect 383580 480 383608 2994
rect 384776 480 384804 3674
rect 384960 3534 384988 64846
rect 385604 62898 385632 65484
rect 386524 63170 386552 65484
rect 387536 64874 387564 65484
rect 387536 64846 387748 64874
rect 386512 63164 386564 63170
rect 386512 63106 386564 63112
rect 387616 63164 387668 63170
rect 387616 63106 387668 63112
rect 385592 62892 385644 62898
rect 385592 62834 385644 62840
rect 386328 62892 386380 62898
rect 386328 62834 386380 62840
rect 386340 5166 386368 62834
rect 386328 5160 386380 5166
rect 386328 5102 386380 5108
rect 387628 3738 387656 63106
rect 387616 3732 387668 3738
rect 387616 3674 387668 3680
rect 384948 3528 385000 3534
rect 384948 3470 385000 3476
rect 387720 3398 387748 64846
rect 388456 63034 388484 65484
rect 388444 63028 388496 63034
rect 388444 62970 388496 62976
rect 389088 63028 389140 63034
rect 389088 62970 389140 62976
rect 389100 5098 389128 62970
rect 389468 62150 389496 65484
rect 390388 64874 390416 65484
rect 390388 64846 390508 64874
rect 389456 62144 389508 62150
rect 389456 62086 389508 62092
rect 390284 62144 390336 62150
rect 390284 62086 390336 62092
rect 389088 5092 389140 5098
rect 389088 5034 389140 5040
rect 390296 4010 390324 62086
rect 389456 4004 389508 4010
rect 389456 3946 389508 3952
rect 390284 4004 390336 4010
rect 390284 3946 390336 3952
rect 388260 3460 388312 3466
rect 388260 3402 388312 3408
rect 385960 3392 386012 3398
rect 385960 3334 386012 3340
rect 387708 3392 387760 3398
rect 387708 3334 387760 3340
rect 385972 480 386000 3334
rect 387156 3120 387208 3126
rect 387156 3062 387208 3068
rect 387168 480 387196 3062
rect 388272 480 388300 3402
rect 389468 480 389496 3946
rect 390480 3466 390508 64846
rect 391400 62490 391428 65484
rect 392320 63374 392348 65484
rect 392308 63368 392360 63374
rect 392308 63310 392360 63316
rect 393228 63368 393280 63374
rect 393228 63310 393280 63316
rect 391388 62484 391440 62490
rect 391388 62426 391440 62432
rect 392584 62484 392636 62490
rect 392584 62426 392636 62432
rect 392596 5030 392624 62426
rect 392584 5024 392636 5030
rect 392584 4966 392636 4972
rect 390652 4140 390704 4146
rect 390652 4082 390704 4088
rect 390468 3460 390520 3466
rect 390468 3402 390520 3408
rect 390664 480 390692 4082
rect 393044 4072 393096 4078
rect 393044 4014 393096 4020
rect 391848 3324 391900 3330
rect 391848 3266 391900 3272
rect 391860 480 391888 3266
rect 393056 480 393084 4014
rect 393240 3330 393268 63310
rect 393332 62354 393360 65484
rect 394252 64874 394280 65484
rect 394252 64846 394556 64874
rect 393320 62348 393372 62354
rect 393320 62290 393372 62296
rect 394528 4962 394556 64846
rect 394608 62348 394660 62354
rect 394608 62290 394660 62296
rect 394516 4956 394568 4962
rect 394516 4898 394568 4904
rect 394620 4078 394648 62290
rect 395264 62150 395292 65484
rect 396184 62354 396212 65484
rect 397196 64874 397224 65484
rect 397196 64846 397316 64874
rect 396172 62348 396224 62354
rect 396172 62290 396224 62296
rect 395252 62144 395304 62150
rect 395252 62086 395304 62092
rect 395988 62144 396040 62150
rect 395988 62086 396040 62092
rect 394608 4072 394660 4078
rect 394608 4014 394660 4020
rect 393228 3324 393280 3330
rect 393228 3266 393280 3272
rect 394240 3256 394292 3262
rect 394240 3198 394292 3204
rect 394252 480 394280 3198
rect 395344 3188 395396 3194
rect 395344 3130 395396 3136
rect 395356 480 395384 3130
rect 396000 3058 396028 62086
rect 397288 4894 397316 64846
rect 398116 62830 398144 65484
rect 398104 62824 398156 62830
rect 398104 62766 398156 62772
rect 398748 62824 398800 62830
rect 398748 62766 398800 62772
rect 397368 62348 397420 62354
rect 397368 62290 397420 62296
rect 397276 4888 397328 4894
rect 397276 4830 397328 4836
rect 397380 4146 397408 62290
rect 397368 4140 397420 4146
rect 397368 4082 397420 4088
rect 398760 3942 398788 62766
rect 399128 62422 399156 65484
rect 399116 62416 399168 62422
rect 399116 62358 399168 62364
rect 400048 4826 400076 65484
rect 400128 62416 400180 62422
rect 400128 62358 400180 62364
rect 398932 4820 398984 4826
rect 398932 4762 398984 4768
rect 400036 4820 400088 4826
rect 400036 4762 400088 4768
rect 397736 3936 397788 3942
rect 397736 3878 397788 3884
rect 398748 3936 398800 3942
rect 398748 3878 398800 3884
rect 396540 3596 396592 3602
rect 396540 3538 396592 3544
rect 395988 3052 396040 3058
rect 395988 2994 396040 3000
rect 396552 480 396580 3538
rect 397748 480 397776 3878
rect 398944 480 398972 4762
rect 400140 3874 400168 62358
rect 401060 62150 401088 65484
rect 401980 62150 402008 65484
rect 402992 62150 403020 65484
rect 403912 64874 403940 65484
rect 403912 64846 404308 64874
rect 401048 62144 401100 62150
rect 401048 62086 401100 62092
rect 401508 62144 401560 62150
rect 401508 62086 401560 62092
rect 401968 62144 402020 62150
rect 401968 62086 402020 62092
rect 402888 62144 402940 62150
rect 402888 62086 402940 62092
rect 402980 62144 403032 62150
rect 402980 62086 403032 62092
rect 404176 62144 404228 62150
rect 404176 62086 404228 62092
rect 400036 3868 400088 3874
rect 400036 3810 400088 3816
rect 400128 3868 400180 3874
rect 400128 3810 400180 3816
rect 400048 1986 400076 3810
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 400048 1958 400168 1986
rect 400140 480 400168 1958
rect 401336 480 401364 3606
rect 401520 3126 401548 62086
rect 402520 5228 402572 5234
rect 402520 5170 402572 5176
rect 401508 3120 401560 3126
rect 401508 3062 401560 3068
rect 402532 480 402560 5170
rect 402900 3670 402928 62086
rect 404188 5302 404216 62086
rect 404176 5296 404228 5302
rect 404176 5238 404228 5244
rect 404280 3806 404308 64846
rect 404924 62898 404952 65484
rect 405844 63170 405872 65484
rect 406856 64874 406884 65484
rect 406856 64846 407068 64874
rect 405832 63164 405884 63170
rect 405832 63106 405884 63112
rect 406936 63164 406988 63170
rect 406936 63106 406988 63112
rect 404912 62892 404964 62898
rect 404912 62834 404964 62840
rect 405648 62892 405700 62898
rect 405648 62834 405700 62840
rect 403624 3800 403676 3806
rect 403624 3742 403676 3748
rect 404268 3800 404320 3806
rect 404268 3742 404320 3748
rect 402888 3664 402940 3670
rect 402888 3606 402940 3612
rect 403636 480 403664 3742
rect 405660 3602 405688 62834
rect 406948 5234 406976 63106
rect 406936 5228 406988 5234
rect 406936 5170 406988 5176
rect 406016 5160 406068 5166
rect 406016 5102 406068 5108
rect 405648 3596 405700 3602
rect 405648 3538 405700 3544
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 404832 480 404860 3470
rect 406028 480 406056 5102
rect 407040 3534 407068 64846
rect 407776 63034 407804 65484
rect 407764 63028 407816 63034
rect 407764 62970 407816 62976
rect 408408 63028 408460 63034
rect 408408 62970 408460 62976
rect 408420 6914 408448 62970
rect 408788 62286 408816 65484
rect 409708 64874 409736 65484
rect 409708 64846 409828 64874
rect 408776 62280 408828 62286
rect 408776 62222 408828 62228
rect 408328 6886 408448 6914
rect 407212 3732 407264 3738
rect 407212 3674 407264 3680
rect 407028 3528 407080 3534
rect 407028 3470 407080 3476
rect 407224 480 407252 3674
rect 408328 3194 408356 6886
rect 409604 5092 409656 5098
rect 409604 5034 409656 5040
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408316 3188 408368 3194
rect 408316 3130 408368 3136
rect 408420 480 408448 3334
rect 409616 480 409644 5034
rect 409800 3398 409828 64846
rect 410524 62280 410576 62286
rect 410524 62222 410576 62228
rect 410536 5370 410564 62222
rect 410720 62150 410748 65484
rect 411640 63374 411668 65484
rect 411628 63368 411680 63374
rect 411628 63310 411680 63316
rect 412548 63368 412600 63374
rect 412548 63310 412600 63316
rect 410708 62144 410760 62150
rect 410708 62086 410760 62092
rect 411168 62144 411220 62150
rect 411168 62086 411220 62092
rect 410524 5364 410576 5370
rect 410524 5306 410576 5312
rect 410800 4004 410852 4010
rect 410800 3946 410852 3952
rect 409788 3392 409840 3398
rect 409788 3334 409840 3340
rect 410812 480 410840 3946
rect 411180 3262 411208 62086
rect 412560 5166 412588 63310
rect 412652 62150 412680 65484
rect 413572 64874 413600 65484
rect 413572 64846 413968 64874
rect 412640 62144 412692 62150
rect 412640 62086 412692 62092
rect 413836 62144 413888 62150
rect 413836 62086 413888 62092
rect 412548 5160 412600 5166
rect 412548 5102 412600 5108
rect 413100 5024 413152 5030
rect 413100 4966 413152 4972
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 411168 3256 411220 3262
rect 411168 3198 411220 3204
rect 411916 480 411944 3402
rect 413112 480 413140 4966
rect 413848 3738 413876 62086
rect 413940 4010 413968 64846
rect 414584 62150 414612 65484
rect 415504 62150 415532 65484
rect 416516 62898 416544 65484
rect 416504 62892 416556 62898
rect 416504 62834 416556 62840
rect 417436 62830 417464 65484
rect 417424 62824 417476 62830
rect 417424 62766 417476 62772
rect 418068 62824 418120 62830
rect 418068 62766 418120 62772
rect 414572 62144 414624 62150
rect 414572 62086 414624 62092
rect 415308 62144 415360 62150
rect 415308 62086 415360 62092
rect 415492 62144 415544 62150
rect 415492 62086 415544 62092
rect 416688 62144 416740 62150
rect 416688 62086 416740 62092
rect 415320 5098 415348 62086
rect 416700 6914 416728 62086
rect 416608 6886 416728 6914
rect 415308 5092 415360 5098
rect 415308 5034 415360 5040
rect 415492 4072 415544 4078
rect 415492 4014 415544 4020
rect 413928 4004 413980 4010
rect 413928 3946 413980 3952
rect 413836 3732 413888 3738
rect 413836 3674 413888 3680
rect 414296 3324 414348 3330
rect 414296 3266 414348 3272
rect 414308 480 414336 3266
rect 415504 480 415532 4014
rect 416608 3330 416636 6886
rect 418080 5030 418108 62766
rect 418448 62422 418476 65484
rect 418436 62416 418488 62422
rect 418436 62358 418488 62364
rect 418068 5024 418120 5030
rect 418068 4966 418120 4972
rect 416688 4956 416740 4962
rect 416688 4898 416740 4904
rect 416596 3324 416648 3330
rect 416596 3266 416648 3272
rect 416700 480 416728 4898
rect 418988 4140 419040 4146
rect 418988 4082 419040 4088
rect 417884 3052 417936 3058
rect 417884 2994 417936 3000
rect 417896 480 417924 2994
rect 419000 480 419028 4082
rect 419368 3466 419396 65484
rect 420380 62422 420408 65484
rect 421300 63034 421328 65484
rect 422312 63102 422340 65484
rect 422300 63096 422352 63102
rect 422300 63038 422352 63044
rect 421288 63028 421340 63034
rect 421288 62970 421340 62976
rect 422208 63028 422260 63034
rect 422208 62970 422260 62976
rect 419448 62416 419500 62422
rect 419448 62358 419500 62364
rect 420368 62416 420420 62422
rect 420368 62358 420420 62364
rect 421564 62416 421616 62422
rect 421564 62358 421616 62364
rect 419460 4146 419488 62358
rect 421576 4962 421604 62358
rect 421564 4956 421616 4962
rect 421564 4898 421616 4904
rect 420184 4888 420236 4894
rect 420184 4830 420236 4836
rect 419448 4140 419500 4146
rect 419448 4082 419500 4088
rect 419356 3460 419408 3466
rect 419356 3402 419408 3408
rect 420196 480 420224 4830
rect 422220 4078 422248 62970
rect 423232 62966 423260 65484
rect 423220 62960 423272 62966
rect 423220 62902 423272 62908
rect 424244 62898 424272 65484
rect 424232 62892 424284 62898
rect 424232 62834 424284 62840
rect 424968 62892 425020 62898
rect 424968 62834 425020 62840
rect 423772 4820 423824 4826
rect 423772 4762 423824 4768
rect 422208 4072 422260 4078
rect 422208 4014 422260 4020
rect 421380 3936 421432 3942
rect 421380 3878 421432 3884
rect 421392 480 421420 3878
rect 422576 3868 422628 3874
rect 422576 3810 422628 3816
rect 422588 480 422616 3810
rect 423784 480 423812 4762
rect 424980 3874 425008 62834
rect 425164 62150 425192 65484
rect 426176 64874 426204 65484
rect 426176 64846 426296 64874
rect 425152 62144 425204 62150
rect 425152 62086 425204 62092
rect 426268 4826 426296 64846
rect 427096 63034 427124 65484
rect 427084 63028 427136 63034
rect 427084 62970 427136 62976
rect 427728 63028 427780 63034
rect 427728 62970 427780 62976
rect 426348 62144 426400 62150
rect 426348 62086 426400 62092
rect 426256 4820 426308 4826
rect 426256 4762 426308 4768
rect 426360 3942 426388 62086
rect 427268 5296 427320 5302
rect 427268 5238 427320 5244
rect 426348 3936 426400 3942
rect 426348 3878 426400 3884
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 426164 3664 426216 3670
rect 426164 3606 426216 3612
rect 424968 3120 425020 3126
rect 424968 3062 425020 3068
rect 424980 480 425008 3062
rect 426176 480 426204 3606
rect 427280 480 427308 5238
rect 427740 3670 427768 62970
rect 428108 62150 428136 65484
rect 428096 62144 428148 62150
rect 428096 62086 428148 62092
rect 429028 4894 429056 65484
rect 430040 62150 430068 65484
rect 430960 62150 430988 65484
rect 431224 62824 431276 62830
rect 431224 62766 431276 62772
rect 429108 62144 429160 62150
rect 429108 62086 429160 62092
rect 430028 62144 430080 62150
rect 430028 62086 430080 62092
rect 430488 62144 430540 62150
rect 430488 62086 430540 62092
rect 430948 62144 431000 62150
rect 430948 62086 431000 62092
rect 429016 4888 429068 4894
rect 429016 4830 429068 4836
rect 428464 3800 428516 3806
rect 428464 3742 428516 3748
rect 427728 3664 427780 3670
rect 427728 3606 427780 3612
rect 428476 480 428504 3742
rect 429120 2854 429148 62086
rect 430500 3806 430528 62086
rect 430856 5228 430908 5234
rect 430856 5170 430908 5176
rect 430488 3800 430540 3806
rect 430488 3742 430540 3748
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 429108 2848 429160 2854
rect 429108 2790 429160 2796
rect 429672 480 429700 3538
rect 430868 480 430896 5170
rect 431236 3058 431264 62766
rect 431972 62150 432000 65484
rect 432892 64874 432920 65484
rect 432892 64846 433288 64874
rect 431868 62144 431920 62150
rect 431868 62086 431920 62092
rect 431960 62144 432012 62150
rect 431960 62086 432012 62092
rect 433156 62144 433208 62150
rect 433156 62086 433208 62092
rect 431224 3052 431276 3058
rect 431224 2994 431276 3000
rect 431880 2922 431908 62086
rect 433168 5302 433196 62086
rect 433156 5296 433208 5302
rect 433156 5238 433208 5244
rect 433260 3602 433288 64846
rect 433904 62218 433932 65484
rect 434824 62966 434852 65484
rect 435836 64874 435864 65484
rect 435836 64846 436048 64874
rect 434812 62960 434864 62966
rect 434812 62902 434864 62908
rect 433892 62212 433944 62218
rect 433892 62154 433944 62160
rect 434444 5364 434496 5370
rect 434444 5306 434496 5312
rect 433248 3596 433300 3602
rect 433248 3538 433300 3544
rect 432052 3528 432104 3534
rect 432052 3470 432104 3476
rect 431868 2916 431920 2922
rect 431868 2858 431920 2864
rect 432064 480 432092 3470
rect 433248 3188 433300 3194
rect 433248 3130 433300 3136
rect 433260 480 433288 3130
rect 434456 480 434484 5306
rect 435548 3392 435600 3398
rect 435548 3334 435600 3340
rect 435560 480 435588 3334
rect 436020 3194 436048 64846
rect 436652 63096 436704 63102
rect 436652 63038 436704 63044
rect 436664 55214 436692 63038
rect 436756 62150 436784 65484
rect 437768 63034 437796 65484
rect 438688 64874 438716 65484
rect 438688 64846 438808 64874
rect 437756 63028 437808 63034
rect 437756 62970 437808 62976
rect 436744 62144 436796 62150
rect 436744 62086 436796 62092
rect 437388 62144 437440 62150
rect 437388 62086 437440 62092
rect 436664 55186 436784 55214
rect 436756 16574 436784 55186
rect 436756 16546 436876 16574
rect 436744 3256 436796 3262
rect 436744 3198 436796 3204
rect 436008 3188 436060 3194
rect 436008 3130 436060 3136
rect 436756 480 436784 3198
rect 436848 2990 436876 16546
rect 437400 3126 437428 62086
rect 437940 5160 437992 5166
rect 437940 5102 437992 5108
rect 437388 3120 437440 3126
rect 437388 3062 437440 3068
rect 436836 2984 436888 2990
rect 436836 2926 436888 2932
rect 437952 480 437980 5102
rect 438780 3534 438808 64846
rect 439700 63238 439728 65484
rect 439688 63232 439740 63238
rect 439688 63174 439740 63180
rect 440148 63232 440200 63238
rect 440148 63174 440200 63180
rect 439504 62212 439556 62218
rect 439504 62154 439556 62160
rect 439516 4010 439544 62154
rect 439504 4004 439556 4010
rect 439504 3946 439556 3952
rect 440160 3738 440188 63174
rect 440620 63170 440648 65484
rect 440608 63164 440660 63170
rect 440608 63106 440660 63112
rect 441528 63164 441580 63170
rect 441528 63106 441580 63112
rect 441436 5092 441488 5098
rect 441436 5034 441488 5040
rect 439136 3732 439188 3738
rect 439136 3674 439188 3680
rect 440148 3732 440200 3738
rect 440148 3674 440200 3680
rect 438768 3528 438820 3534
rect 438768 3470 438820 3476
rect 439148 480 439176 3674
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440344 480 440372 3334
rect 441448 2530 441476 5034
rect 441540 3398 441568 63106
rect 441632 62422 441660 65484
rect 442552 62830 442580 65484
rect 442540 62824 442592 62830
rect 442540 62766 442592 62772
rect 441620 62416 441672 62422
rect 441620 62358 441672 62364
rect 442908 62416 442960 62422
rect 442908 62358 442960 62364
rect 442920 4214 442948 62358
rect 443564 62150 443592 65484
rect 444484 63102 444512 65484
rect 445496 63374 445524 65484
rect 445484 63368 445536 63374
rect 445484 63310 445536 63316
rect 444472 63096 444524 63102
rect 444472 63038 444524 63044
rect 446312 62892 446364 62898
rect 446312 62834 446364 62840
rect 443552 62144 443604 62150
rect 443552 62086 443604 62092
rect 444288 62144 444340 62150
rect 444288 62086 444340 62092
rect 442908 4208 442960 4214
rect 442908 4150 442960 4156
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 444300 3330 444328 62086
rect 446324 55214 446352 62834
rect 446416 62150 446444 65484
rect 447428 62150 447456 65484
rect 448348 64874 448376 65484
rect 448348 64846 448468 64874
rect 446404 62144 446456 62150
rect 446404 62086 446456 62092
rect 447048 62144 447100 62150
rect 447048 62086 447100 62092
rect 447416 62144 447468 62150
rect 447416 62086 447468 62092
rect 448244 62144 448296 62150
rect 448244 62086 448296 62092
rect 446324 55186 446444 55214
rect 445024 5024 445076 5030
rect 445024 4966 445076 4972
rect 442632 3324 442684 3330
rect 442632 3266 442684 3272
rect 444288 3324 444340 3330
rect 444288 3266 444340 3272
rect 441448 2502 441568 2530
rect 441540 480 441568 2502
rect 442644 480 442672 3266
rect 443828 3052 443880 3058
rect 443828 2994 443880 3000
rect 443840 480 443868 2994
rect 445036 480 445064 4966
rect 446416 4418 446444 55186
rect 447060 5234 447088 62086
rect 447048 5228 447100 5234
rect 447048 5170 447100 5176
rect 446404 4412 446456 4418
rect 446404 4354 446456 4360
rect 446220 4140 446272 4146
rect 446220 4082 446272 4088
rect 446232 480 446260 4082
rect 448256 3466 448284 62086
rect 447416 3460 447468 3466
rect 447416 3402 447468 3408
rect 448244 3460 448296 3466
rect 448244 3402 448296 3408
rect 447428 480 447456 3402
rect 448440 3330 448468 64846
rect 449164 63368 449216 63374
rect 449164 63310 449216 63316
rect 448612 4956 448664 4962
rect 448612 4898 448664 4904
rect 448428 3324 448480 3330
rect 448428 3266 448480 3272
rect 448624 480 448652 4898
rect 449176 3058 449204 63310
rect 449360 62150 449388 65484
rect 450280 62286 450308 65484
rect 451292 63170 451320 65484
rect 451280 63164 451332 63170
rect 451280 63106 451332 63112
rect 452212 62626 452240 65484
rect 452200 62620 452252 62626
rect 452200 62562 452252 62568
rect 450268 62280 450320 62286
rect 450268 62222 450320 62228
rect 451188 62280 451240 62286
rect 451188 62222 451240 62228
rect 449348 62144 449400 62150
rect 449348 62086 449400 62092
rect 449808 62144 449860 62150
rect 449808 62086 449860 62092
rect 449820 5098 449848 62086
rect 449808 5092 449860 5098
rect 449808 5034 449860 5040
rect 451200 4146 451228 62222
rect 453224 62150 453252 65484
rect 454144 63306 454172 65484
rect 455156 64874 455184 65484
rect 455156 64846 455368 64874
rect 454132 63300 454184 63306
rect 454132 63242 454184 63248
rect 454684 63028 454736 63034
rect 454684 62970 454736 62976
rect 453304 62620 453356 62626
rect 453304 62562 453356 62568
rect 453212 62144 453264 62150
rect 453212 62086 453264 62092
rect 453316 5166 453344 62562
rect 453948 62144 454000 62150
rect 453948 62086 454000 62092
rect 453304 5160 453356 5166
rect 453304 5102 453356 5108
rect 452108 4412 452160 4418
rect 452108 4354 452160 4360
rect 451188 4140 451240 4146
rect 451188 4082 451240 4088
rect 449808 4072 449860 4078
rect 449808 4014 449860 4020
rect 449164 3052 449216 3058
rect 449164 2994 449216 3000
rect 449820 480 449848 4014
rect 450912 2984 450964 2990
rect 450912 2926 450964 2932
rect 450924 480 450952 2926
rect 452120 480 452148 4354
rect 453960 4010 453988 62086
rect 454696 5370 454724 62970
rect 454684 5364 454736 5370
rect 454684 5306 454736 5312
rect 455340 5030 455368 64846
rect 456076 62150 456104 65484
rect 457088 63374 457116 65484
rect 458008 64874 458036 65484
rect 458008 64846 458128 64874
rect 457076 63368 457128 63374
rect 457076 63310 457128 63316
rect 456064 62144 456116 62150
rect 456064 62086 456116 62092
rect 456708 62144 456760 62150
rect 456708 62086 456760 62092
rect 455328 5024 455380 5030
rect 455328 4966 455380 4972
rect 455696 4820 455748 4826
rect 455696 4762 455748 4768
rect 453948 4004 454000 4010
rect 453948 3946 454000 3952
rect 453304 3868 453356 3874
rect 453304 3810 453356 3816
rect 453316 480 453344 3810
rect 454500 3800 454552 3806
rect 454500 3742 454552 3748
rect 454512 480 454540 3742
rect 455708 480 455736 4762
rect 456720 4078 456748 62086
rect 458100 4962 458128 64846
rect 459020 62150 459048 65484
rect 459940 62150 459968 65484
rect 460952 62150 460980 65484
rect 461872 64874 461900 65484
rect 461872 64846 462268 64874
rect 459008 62144 459060 62150
rect 459008 62086 459060 62092
rect 459468 62144 459520 62150
rect 459468 62086 459520 62092
rect 459928 62144 459980 62150
rect 459928 62086 459980 62092
rect 460848 62144 460900 62150
rect 460848 62086 460900 62092
rect 460940 62144 460992 62150
rect 460940 62086 460992 62092
rect 462136 62144 462188 62150
rect 462136 62086 462188 62092
rect 458088 4956 458140 4962
rect 458088 4898 458140 4904
rect 459192 4888 459244 4894
rect 459192 4830 459244 4836
rect 456708 4072 456760 4078
rect 456708 4014 456760 4020
rect 456892 3664 456944 3670
rect 456892 3606 456944 3612
rect 456904 480 456932 3606
rect 458088 2848 458140 2854
rect 458088 2790 458140 2796
rect 458100 480 458128 2790
rect 459204 480 459232 4830
rect 459480 3670 459508 62086
rect 460860 3874 460888 62086
rect 462148 4894 462176 62086
rect 462136 4888 462188 4894
rect 462136 4830 462188 4836
rect 460388 3868 460440 3874
rect 460388 3810 460440 3816
rect 460848 3868 460900 3874
rect 460848 3810 460900 3816
rect 459468 3664 459520 3670
rect 459468 3606 459520 3612
rect 460400 480 460428 3810
rect 462240 3754 462268 64846
rect 462884 63238 462912 65484
rect 462872 63232 462924 63238
rect 462872 63174 462924 63180
rect 463804 63034 463832 65484
rect 464344 63096 464396 63102
rect 464344 63038 464396 63044
rect 463792 63028 463844 63034
rect 463792 62970 463844 62976
rect 462780 5296 462832 5302
rect 462780 5238 462832 5244
rect 462240 3726 462452 3754
rect 462424 3670 462452 3726
rect 462412 3664 462464 3670
rect 462412 3606 462464 3612
rect 461584 2916 461636 2922
rect 461584 2858 461636 2864
rect 461596 480 461624 2858
rect 462792 480 462820 5238
rect 463976 3596 464028 3602
rect 463976 3538 464028 3544
rect 463988 480 464016 3538
rect 464356 2922 464384 63038
rect 464816 62898 464844 65484
rect 465172 62960 465224 62966
rect 465172 62902 465224 62908
rect 464804 62892 464856 62898
rect 464804 62834 464856 62840
rect 465184 16574 465212 62902
rect 465736 62150 465764 65484
rect 466748 62150 466776 65484
rect 467668 63170 467696 65484
rect 468484 63300 468536 63306
rect 468484 63242 468536 63248
rect 467104 63164 467156 63170
rect 467104 63106 467156 63112
rect 467656 63164 467708 63170
rect 467656 63106 467708 63112
rect 465724 62144 465776 62150
rect 465724 62086 465776 62092
rect 466368 62144 466420 62150
rect 466368 62086 466420 62092
rect 466736 62144 466788 62150
rect 466736 62086 466788 62092
rect 465184 16546 466316 16574
rect 465172 3936 465224 3942
rect 465172 3878 465224 3884
rect 464344 2916 464396 2922
rect 464344 2858 464396 2864
rect 465184 480 465212 3878
rect 466288 480 466316 16546
rect 466380 3738 466408 62086
rect 466368 3732 466420 3738
rect 466368 3674 466420 3680
rect 467116 3602 467144 63106
rect 467748 62144 467800 62150
rect 467748 62086 467800 62092
rect 467760 4826 467788 62086
rect 467748 4820 467800 4826
rect 467748 4762 467800 4768
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 467564 3596 467616 3602
rect 467564 3538 467616 3544
rect 467576 3194 467604 3538
rect 467472 3188 467524 3194
rect 467472 3130 467524 3136
rect 467564 3188 467616 3194
rect 467564 3130 467616 3136
rect 467484 480 467512 3130
rect 468496 2854 468524 63242
rect 468680 62966 468708 65484
rect 468668 62960 468720 62966
rect 468668 62902 468720 62908
rect 469600 62218 469628 65484
rect 470612 63442 470640 65484
rect 471532 64874 471560 65484
rect 471532 64846 471928 64874
rect 470600 63436 470652 63442
rect 470600 63378 470652 63384
rect 471244 63368 471296 63374
rect 471244 63310 471296 63316
rect 469588 62212 469640 62218
rect 469588 62154 469640 62160
rect 469864 5364 469916 5370
rect 469864 5306 469916 5312
rect 468668 3120 468720 3126
rect 468668 3062 468720 3068
rect 468484 2848 468536 2854
rect 468484 2790 468536 2796
rect 468680 480 468708 3062
rect 469876 480 469904 5306
rect 471060 3528 471112 3534
rect 471060 3470 471112 3476
rect 471072 480 471100 3470
rect 471256 2922 471284 63310
rect 471900 3534 471928 64846
rect 472544 62150 472572 65484
rect 473464 62218 473492 65484
rect 474476 63102 474504 65484
rect 474464 63096 474516 63102
rect 474464 63038 474516 63044
rect 474004 62824 474056 62830
rect 474004 62766 474056 62772
rect 472624 62212 472676 62218
rect 472624 62154 472676 62160
rect 473452 62212 473504 62218
rect 473452 62154 473504 62160
rect 472532 62144 472584 62150
rect 472532 62086 472584 62092
rect 472636 5506 472664 62154
rect 473268 62144 473320 62150
rect 473268 62086 473320 62092
rect 473280 6186 473308 62086
rect 473268 6180 473320 6186
rect 473268 6122 473320 6128
rect 472624 5500 472676 5506
rect 472624 5442 472676 5448
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 471888 3528 471940 3534
rect 471888 3470 471940 3476
rect 471244 2916 471296 2922
rect 471244 2858 471296 2864
rect 472268 480 472296 3538
rect 474016 3534 474044 62766
rect 475396 62150 475424 65484
rect 476408 62490 476436 65484
rect 477328 62626 477356 65484
rect 477316 62620 477368 62626
rect 477316 62562 477368 62568
rect 478340 62558 478368 65484
rect 478328 62552 478380 62558
rect 478328 62494 478380 62500
rect 476396 62484 476448 62490
rect 476396 62426 476448 62432
rect 476764 62212 476816 62218
rect 476764 62154 476816 62160
rect 475384 62144 475436 62150
rect 475384 62086 475436 62092
rect 476028 62144 476080 62150
rect 476028 62086 476080 62092
rect 476040 5370 476068 62086
rect 476028 5364 476080 5370
rect 476028 5306 476080 5312
rect 476776 3738 476804 62154
rect 479260 62150 479288 65484
rect 479524 62552 479576 62558
rect 479524 62494 479576 62500
rect 479248 62144 479300 62150
rect 479248 62086 479300 62092
rect 479536 8974 479564 62494
rect 480272 62218 480300 65484
rect 481192 62286 481220 65484
rect 482204 63306 482232 65484
rect 482192 63300 482244 63306
rect 482192 63242 482244 63248
rect 482928 63300 482980 63306
rect 482928 63242 482980 63248
rect 482284 63232 482336 63238
rect 482284 63174 482336 63180
rect 481180 62280 481232 62286
rect 481180 62222 481232 62228
rect 480260 62212 480312 62218
rect 480260 62154 480312 62160
rect 480168 62144 480220 62150
rect 480168 62086 480220 62092
rect 479524 8968 479576 8974
rect 479524 8910 479576 8916
rect 476764 3732 476816 3738
rect 476764 3674 476816 3680
rect 480180 3534 480208 62086
rect 480536 5228 480588 5234
rect 480536 5170 480588 5176
rect 474004 3528 474056 3534
rect 474004 3470 474056 3476
rect 475752 3528 475804 3534
rect 475752 3470 475804 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 473452 3392 473504 3398
rect 473452 3334 473504 3340
rect 473464 480 473492 3334
rect 474556 3052 474608 3058
rect 474556 2994 474608 3000
rect 474568 480 474596 2994
rect 475764 480 475792 3470
rect 476948 3256 477000 3262
rect 476948 3198 477000 3204
rect 476960 480 476988 3198
rect 478144 3120 478196 3126
rect 478144 3062 478196 3068
rect 478156 480 478184 3062
rect 479340 2984 479392 2990
rect 479340 2926 479392 2932
rect 479352 480 479380 2926
rect 480548 480 480576 5170
rect 481732 3460 481784 3466
rect 481732 3402 481784 3408
rect 481744 480 481772 3402
rect 482296 3330 482324 63174
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482284 3324 482336 3330
rect 482284 3266 482336 3272
rect 482848 480 482876 3334
rect 482940 2990 482968 63242
rect 483124 62422 483152 65484
rect 484136 64874 484164 65484
rect 484136 64846 484348 64874
rect 483112 62416 483164 62422
rect 483112 62358 483164 62364
rect 483664 62212 483716 62218
rect 483664 62154 483716 62160
rect 483676 3126 483704 62154
rect 484320 5302 484348 64846
rect 485056 62150 485084 65484
rect 486068 62762 486096 65484
rect 486988 64874 487016 65484
rect 486988 64846 487108 64874
rect 486056 62756 486108 62762
rect 486056 62698 486108 62704
rect 485136 62280 485188 62286
rect 485136 62222 485188 62228
rect 485044 62144 485096 62150
rect 485044 62086 485096 62092
rect 485148 5438 485176 62222
rect 485688 62144 485740 62150
rect 485688 62086 485740 62092
rect 485136 5432 485188 5438
rect 485136 5374 485188 5380
rect 484308 5296 484360 5302
rect 484308 5238 484360 5244
rect 484032 5092 484084 5098
rect 484032 5034 484084 5040
rect 483664 3120 483716 3126
rect 483664 3062 483716 3068
rect 482928 2984 482980 2990
rect 482928 2926 482980 2932
rect 484044 480 484072 5034
rect 485228 4140 485280 4146
rect 485228 4082 485280 4088
rect 485240 480 485268 4082
rect 485700 3466 485728 62086
rect 487080 5098 487108 64846
rect 487804 62960 487856 62966
rect 487804 62902 487856 62908
rect 487620 5160 487672 5166
rect 487620 5102 487672 5108
rect 487068 5092 487120 5098
rect 487068 5034 487120 5040
rect 485688 3460 485740 3466
rect 485688 3402 485740 3408
rect 486424 3188 486476 3194
rect 486424 3130 486476 3136
rect 486436 480 486464 3130
rect 487632 480 487660 5102
rect 487816 4146 487844 62902
rect 488000 62694 488028 65484
rect 487988 62688 488040 62694
rect 487988 62630 488040 62636
rect 488920 62150 488948 65484
rect 489932 63238 489960 65484
rect 489920 63232 489972 63238
rect 489920 63174 489972 63180
rect 490852 63102 490880 65484
rect 490564 63096 490616 63102
rect 490564 63038 490616 63044
rect 490840 63096 490892 63102
rect 490840 63038 490892 63044
rect 488908 62144 488960 62150
rect 488908 62086 488960 62092
rect 489828 62144 489880 62150
rect 489828 62086 489880 62092
rect 487804 4140 487856 4146
rect 487804 4082 487856 4088
rect 488816 4004 488868 4010
rect 488816 3946 488868 3952
rect 488828 480 488856 3946
rect 489840 3262 489868 62086
rect 489828 3256 489880 3262
rect 489828 3198 489880 3204
rect 490576 3058 490604 63038
rect 491864 62966 491892 65484
rect 491852 62960 491904 62966
rect 491852 62902 491904 62908
rect 492784 62898 492812 65484
rect 493796 63306 493824 65484
rect 494716 63374 494744 65484
rect 494704 63368 494756 63374
rect 494704 63310 494756 63316
rect 495348 63368 495400 63374
rect 495348 63310 495400 63316
rect 493784 63300 493836 63306
rect 493784 63242 493836 63248
rect 492772 62892 492824 62898
rect 492772 62834 492824 62840
rect 493968 62892 494020 62898
rect 493968 62834 494020 62840
rect 493980 5166 494008 62834
rect 493968 5160 494020 5166
rect 493968 5102 494020 5108
rect 491116 5024 491168 5030
rect 491116 4966 491168 4972
rect 490564 3052 490616 3058
rect 490564 2994 490616 3000
rect 489920 2848 489972 2854
rect 489920 2790 489972 2796
rect 489932 480 489960 2790
rect 491128 480 491156 4966
rect 494704 4956 494756 4962
rect 494704 4898 494756 4904
rect 492312 4072 492364 4078
rect 492312 4014 492364 4020
rect 492324 480 492352 4014
rect 493508 2916 493560 2922
rect 493508 2858 493560 2864
rect 493520 480 493548 2858
rect 494716 480 494744 4898
rect 495360 3398 495388 63310
rect 495728 62150 495756 65484
rect 496648 63306 496676 65484
rect 496636 63300 496688 63306
rect 496636 63242 496688 63248
rect 497660 62898 497688 65484
rect 497648 62892 497700 62898
rect 497648 62834 497700 62840
rect 497464 62824 497516 62830
rect 497464 62766 497516 62772
rect 495716 62144 495768 62150
rect 495716 62086 495768 62092
rect 497096 3936 497148 3942
rect 497096 3878 497148 3884
rect 495900 3868 495952 3874
rect 495900 3810 495952 3816
rect 495348 3392 495400 3398
rect 495348 3334 495400 3340
rect 495912 480 495940 3810
rect 497108 480 497136 3878
rect 497476 3874 497504 62766
rect 498580 62150 498608 65484
rect 499592 63510 499620 65484
rect 499580 63504 499632 63510
rect 499580 63446 499632 63452
rect 500512 63034 500540 65484
rect 500316 63028 500368 63034
rect 500316 62970 500368 62976
rect 500500 63028 500552 63034
rect 500500 62970 500552 62976
rect 497556 62144 497608 62150
rect 497556 62086 497608 62092
rect 498568 62144 498620 62150
rect 498568 62086 498620 62092
rect 500224 62144 500276 62150
rect 500224 62086 500276 62092
rect 497568 5234 497596 62086
rect 497556 5228 497608 5234
rect 497556 5170 497608 5176
rect 500236 5030 500264 62086
rect 500224 5024 500276 5030
rect 500224 4966 500276 4972
rect 498200 4888 498252 4894
rect 498200 4830 498252 4836
rect 497464 3868 497516 3874
rect 497464 3810 497516 3816
rect 498212 480 498240 4830
rect 500328 4214 500356 62970
rect 501524 62150 501552 65484
rect 502444 62150 502472 65484
rect 503456 63170 503484 65484
rect 502984 63164 503036 63170
rect 502984 63106 503036 63112
rect 503444 63164 503496 63170
rect 503444 63106 503496 63112
rect 501512 62144 501564 62150
rect 501512 62086 501564 62092
rect 502248 62144 502300 62150
rect 502248 62086 502300 62092
rect 502432 62144 502484 62150
rect 502432 62086 502484 62092
rect 502260 4894 502288 62086
rect 502248 4888 502300 4894
rect 502248 4830 502300 4836
rect 500316 4208 500368 4214
rect 500316 4150 500368 4156
rect 501788 4208 501840 4214
rect 501788 4150 501840 4156
rect 499396 3800 499448 3806
rect 499396 3742 499448 3748
rect 499408 480 499436 3742
rect 500592 3324 500644 3330
rect 500592 3266 500644 3272
rect 500604 480 500632 3266
rect 501800 480 501828 4150
rect 502892 3868 502944 3874
rect 502892 3810 502944 3816
rect 502904 1986 502932 3810
rect 502996 3670 503024 63106
rect 504376 62150 504404 65484
rect 505388 62490 505416 65484
rect 506308 63238 506336 65484
rect 506296 63232 506348 63238
rect 506296 63174 506348 63180
rect 505376 62484 505428 62490
rect 505376 62426 505428 62432
rect 507320 62150 507348 65484
rect 508240 62150 508268 65484
rect 509252 63442 509280 65484
rect 508504 63436 508556 63442
rect 508504 63378 508556 63384
rect 509240 63436 509292 63442
rect 509240 63378 509292 63384
rect 503628 62144 503680 62150
rect 503628 62086 503680 62092
rect 504364 62144 504416 62150
rect 504364 62086 504416 62092
rect 505008 62144 505060 62150
rect 505008 62086 505060 62092
rect 507308 62144 507360 62150
rect 507308 62086 507360 62092
rect 507768 62144 507820 62150
rect 507768 62086 507820 62092
rect 508228 62144 508280 62150
rect 508228 62086 508280 62092
rect 502984 3664 503036 3670
rect 502984 3606 503036 3612
rect 503640 3194 503668 62086
rect 505020 4962 505048 62086
rect 505008 4956 505060 4962
rect 505008 4898 505060 4904
rect 507780 4826 507808 62086
rect 505376 4820 505428 4826
rect 505376 4762 505428 4768
rect 507768 4820 507820 4826
rect 507768 4762 507820 4768
rect 504180 3324 504232 3330
rect 504180 3266 504232 3272
rect 503628 3188 503680 3194
rect 503628 3130 503680 3136
rect 502904 1958 503024 1986
rect 502996 480 503024 1958
rect 504192 480 504220 3266
rect 505388 480 505416 4762
rect 507676 4140 507728 4146
rect 507676 4082 507728 4088
rect 506480 3664 506532 3670
rect 506480 3606 506532 3612
rect 506492 480 506520 3606
rect 507688 480 507716 4082
rect 508516 3330 508544 63378
rect 510172 62218 510200 65484
rect 510160 62212 510212 62218
rect 510160 62154 510212 62160
rect 511184 62150 511212 65484
rect 511264 62212 511316 62218
rect 511264 62154 511316 62160
rect 509148 62144 509200 62150
rect 509148 62086 509200 62092
rect 511172 62144 511224 62150
rect 511172 62086 511224 62092
rect 508872 5500 508924 5506
rect 508872 5442 508924 5448
rect 508504 3324 508556 3330
rect 508504 3266 508556 3272
rect 508884 480 508912 5442
rect 509160 4078 509188 62086
rect 511276 32434 511304 62154
rect 512104 62150 512132 65484
rect 511908 62144 511960 62150
rect 511908 62086 511960 62092
rect 512092 62144 512144 62150
rect 512092 62086 512144 62092
rect 511264 32428 511316 32434
rect 511264 32370 511316 32376
rect 511920 4146 511948 62086
rect 513116 61470 513144 65484
rect 513932 62552 513984 62558
rect 513932 62494 513984 62500
rect 513196 62144 513248 62150
rect 513196 62086 513248 62092
rect 513104 61464 513156 61470
rect 513104 61406 513156 61412
rect 512460 6180 512512 6186
rect 512460 6122 512512 6128
rect 511908 4140 511960 4146
rect 511908 4082 511960 4088
rect 509148 4072 509200 4078
rect 509148 4014 509200 4020
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 510068 3324 510120 3330
rect 510068 3266 510120 3272
rect 510080 480 510108 3266
rect 511276 480 511304 3538
rect 512472 480 512500 6122
rect 513208 4010 513236 62086
rect 513944 55214 513972 62494
rect 514036 62150 514064 65484
rect 515048 62150 515076 65484
rect 515968 62626 515996 65484
rect 515496 62620 515548 62626
rect 515496 62562 515548 62568
rect 515956 62620 516008 62626
rect 515956 62562 516008 62568
rect 515404 62416 515456 62422
rect 515404 62358 515456 62364
rect 514024 62144 514076 62150
rect 514024 62086 514076 62092
rect 514668 62144 514720 62150
rect 514668 62086 514720 62092
rect 515036 62144 515088 62150
rect 515036 62086 515088 62092
rect 513944 55186 514064 55214
rect 513196 4004 513248 4010
rect 513196 3946 513248 3952
rect 513564 3732 513616 3738
rect 513564 3674 513616 3680
rect 513576 480 513604 3674
rect 514036 3602 514064 55186
rect 514680 3942 514708 62086
rect 514668 3936 514720 3942
rect 514668 3878 514720 3884
rect 514024 3596 514076 3602
rect 514024 3538 514076 3544
rect 514760 3052 514812 3058
rect 514760 2994 514812 3000
rect 514772 480 514800 2994
rect 515416 2922 515444 62358
rect 515508 3058 515536 62562
rect 516980 62150 517008 65484
rect 517520 62620 517572 62626
rect 517520 62562 517572 62568
rect 516048 62144 516100 62150
rect 516048 62086 516100 62092
rect 516968 62144 517020 62150
rect 516968 62086 517020 62092
rect 517428 62144 517480 62150
rect 517428 62086 517480 62092
rect 515956 5364 516008 5370
rect 515956 5306 516008 5312
rect 515496 3052 515548 3058
rect 515496 2994 515548 3000
rect 515404 2916 515456 2922
rect 515404 2858 515456 2864
rect 515968 480 515996 5306
rect 516060 3874 516088 62086
rect 516048 3868 516100 3874
rect 516048 3810 516100 3816
rect 517440 3738 517468 62086
rect 517532 61538 517560 62562
rect 517900 62150 517928 65484
rect 518912 62150 518940 65484
rect 519832 62558 519860 65484
rect 519820 62552 519872 62558
rect 519820 62494 519872 62500
rect 520844 62150 520872 65484
rect 517888 62144 517940 62150
rect 517888 62086 517940 62092
rect 518808 62144 518860 62150
rect 518808 62086 518860 62092
rect 518900 62144 518952 62150
rect 518900 62086 518952 62092
rect 520188 62144 520240 62150
rect 520188 62086 520240 62092
rect 520832 62144 520884 62150
rect 520832 62086 520884 62092
rect 521568 62144 521620 62150
rect 521568 62086 521620 62092
rect 517520 61532 517572 61538
rect 517520 61474 517572 61480
rect 518820 3806 518848 62086
rect 520200 8974 520228 62086
rect 519544 8968 519596 8974
rect 519544 8910 519596 8916
rect 520188 8968 520240 8974
rect 520188 8910 520240 8916
rect 518808 3800 518860 3806
rect 518808 3742 518860 3748
rect 517428 3732 517480 3738
rect 517428 3674 517480 3680
rect 517152 3596 517204 3602
rect 517152 3538 517204 3544
rect 517164 480 517192 3538
rect 518348 3052 518400 3058
rect 518348 2994 518400 3000
rect 518360 480 518388 2994
rect 519556 480 519584 8910
rect 521580 3670 521608 62086
rect 521764 61402 521792 65484
rect 522776 64874 522804 65484
rect 522776 64846 522896 64874
rect 521752 61396 521804 61402
rect 521752 61338 521804 61344
rect 521568 3664 521620 3670
rect 521568 3606 521620 3612
rect 520740 3528 520792 3534
rect 520740 3470 520792 3476
rect 520752 480 520780 3470
rect 522868 3194 522896 64846
rect 523696 62626 523724 65484
rect 523684 62620 523736 62626
rect 523684 62562 523736 62568
rect 524708 62354 524736 65484
rect 525064 62756 525116 62762
rect 525064 62698 525116 62704
rect 524696 62348 524748 62354
rect 524696 62290 524748 62296
rect 523040 5432 523092 5438
rect 523040 5374 523092 5380
rect 522856 3188 522908 3194
rect 522856 3130 522908 3136
rect 521844 3120 521896 3126
rect 521844 3062 521896 3068
rect 521856 480 521884 3062
rect 523052 480 523080 5374
rect 525076 3602 525104 62698
rect 525628 62422 525656 65484
rect 526444 62688 526496 62694
rect 526444 62630 526496 62636
rect 525616 62416 525668 62422
rect 525616 62358 525668 62364
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 526456 3126 526484 62630
rect 526640 62150 526668 65484
rect 527560 62150 527588 65484
rect 528572 62762 528600 65484
rect 529492 62830 529520 65484
rect 532056 63096 532108 63102
rect 532056 63038 532108 63044
rect 529204 62824 529256 62830
rect 529204 62766 529256 62772
rect 529480 62824 529532 62830
rect 529480 62766 529532 62772
rect 528560 62756 528612 62762
rect 528560 62698 528612 62704
rect 526628 62144 526680 62150
rect 526628 62086 526680 62092
rect 527088 62144 527140 62150
rect 527088 62086 527140 62092
rect 527548 62144 527600 62150
rect 527548 62086 527600 62092
rect 528468 62144 528520 62150
rect 528468 62086 528520 62092
rect 526628 5296 526680 5302
rect 526628 5238 526680 5244
rect 526444 3120 526496 3126
rect 526444 3062 526496 3068
rect 525432 3052 525484 3058
rect 525432 2994 525484 3000
rect 524236 2984 524288 2990
rect 524236 2926 524288 2932
rect 524248 480 524276 2926
rect 525444 480 525472 2994
rect 526640 480 526668 5238
rect 527100 3534 527128 62086
rect 527088 3528 527140 3534
rect 527088 3470 527140 3476
rect 528480 3466 528508 62086
rect 529216 4214 529244 62766
rect 531964 62348 532016 62354
rect 531964 62290 532016 62296
rect 530124 5092 530176 5098
rect 530124 5034 530176 5040
rect 529204 4208 529256 4214
rect 529204 4150 529256 4156
rect 529020 3596 529072 3602
rect 529020 3538 529072 3544
rect 527824 3460 527876 3466
rect 527824 3402 527876 3408
rect 528468 3460 528520 3466
rect 528468 3402 528520 3408
rect 527836 480 527864 3402
rect 529032 480 529060 3538
rect 530136 480 530164 5034
rect 531976 3126 532004 62290
rect 532068 3602 532096 63038
rect 533356 60722 533384 637735
rect 533448 458182 533476 640018
rect 536116 471986 536144 641446
rect 569316 641436 569368 641442
rect 569316 641378 569368 641384
rect 558276 641368 558328 641374
rect 558276 641310 558328 641316
rect 551376 641164 551428 641170
rect 551376 641106 551428 641112
rect 547236 640756 547288 640762
rect 547236 640698 547288 640704
rect 543004 640620 543056 640626
rect 543004 640562 543056 640568
rect 538956 640280 539008 640286
rect 538956 640222 539008 640228
rect 537576 640212 537628 640218
rect 537576 640154 537628 640160
rect 536196 640144 536248 640150
rect 536196 640086 536248 640092
rect 536208 511970 536236 640086
rect 537484 638580 537536 638586
rect 537484 638522 537536 638528
rect 536196 511964 536248 511970
rect 536196 511906 536248 511912
rect 536104 471980 536156 471986
rect 536104 471922 536156 471928
rect 533436 458176 533488 458182
rect 533436 458118 533488 458124
rect 537496 379506 537524 638522
rect 537588 564398 537616 640154
rect 538864 638376 538916 638382
rect 538864 638318 538916 638324
rect 537576 564392 537628 564398
rect 537576 564334 537628 564340
rect 537484 379500 537536 379506
rect 537484 379442 537536 379448
rect 538876 273222 538904 638318
rect 538968 618254 538996 640222
rect 540244 638988 540296 638994
rect 540244 638930 540296 638936
rect 538956 618248 539008 618254
rect 538956 618190 539008 618196
rect 538864 273216 538916 273222
rect 538864 273158 538916 273164
rect 540256 86970 540284 638930
rect 543016 206990 543044 640562
rect 544476 639532 544528 639538
rect 544476 639474 544528 639480
rect 544384 638172 544436 638178
rect 544384 638114 544436 638120
rect 544396 219434 544424 638114
rect 544488 245614 544516 639474
rect 547144 638104 547196 638110
rect 547144 638046 547196 638052
rect 544476 245608 544528 245614
rect 544476 245550 544528 245556
rect 544384 219428 544436 219434
rect 544384 219370 544436 219376
rect 543004 206984 543056 206990
rect 543004 206926 543056 206932
rect 547156 179382 547184 638046
rect 547248 299470 547276 640698
rect 548616 639736 548668 639742
rect 548616 639678 548668 639684
rect 548524 638036 548576 638042
rect 548524 637978 548576 637984
rect 547236 299464 547288 299470
rect 547236 299406 547288 299412
rect 547144 179376 547196 179382
rect 547144 179318 547196 179324
rect 548536 139398 548564 637978
rect 548628 353258 548656 639678
rect 551284 637900 551336 637906
rect 551284 637842 551336 637848
rect 548616 353252 548668 353258
rect 548616 353194 548668 353200
rect 548524 139392 548576 139398
rect 548524 139334 548576 139340
rect 551296 100706 551324 637842
rect 551388 405686 551416 641106
rect 556802 639296 556858 639305
rect 556802 639231 556858 639240
rect 555422 639024 555478 639033
rect 555422 638959 555478 638968
rect 551376 405680 551428 405686
rect 551376 405622 551428 405628
rect 551284 100700 551336 100706
rect 551284 100642 551336 100648
rect 540244 86964 540296 86970
rect 540244 86906 540296 86912
rect 538864 63504 538916 63510
rect 538864 63446 538916 63452
rect 533436 63368 533488 63374
rect 533436 63310 533488 63316
rect 533344 60716 533396 60722
rect 533344 60658 533396 60664
rect 532056 3596 532108 3602
rect 532056 3538 532108 3544
rect 533448 3262 533476 63310
rect 537484 63300 537536 63306
rect 537484 63242 537536 63248
rect 535460 62960 535512 62966
rect 535460 62902 535512 62908
rect 534724 62552 534776 62558
rect 534724 62494 534776 62500
rect 533712 4208 533764 4214
rect 533712 4150 533764 4156
rect 532516 3256 532568 3262
rect 532516 3198 532568 3204
rect 533436 3256 533488 3262
rect 533436 3198 533488 3204
rect 531320 3120 531372 3126
rect 531320 3062 531372 3068
rect 531964 3120 532016 3126
rect 531964 3062 532016 3068
rect 531332 480 531360 3062
rect 532528 480 532556 3198
rect 533724 480 533752 4150
rect 534736 3058 534764 62494
rect 535472 16574 535500 62902
rect 535472 16546 536144 16574
rect 534908 3596 534960 3602
rect 534908 3538 534960 3544
rect 534724 3052 534776 3058
rect 534724 2994 534776 3000
rect 534920 480 534948 3538
rect 536116 480 536144 16546
rect 537208 5160 537260 5166
rect 537208 5102 537260 5108
rect 537220 480 537248 5102
rect 537496 2990 537524 63242
rect 538404 3256 538456 3262
rect 538404 3198 538456 3204
rect 537484 2984 537536 2990
rect 537484 2926 537536 2932
rect 538416 480 538444 3198
rect 538876 2854 538904 63446
rect 548524 63436 548576 63442
rect 548524 63378 548576 63384
rect 547144 63232 547196 63238
rect 547144 63174 547196 63180
rect 544384 63164 544436 63170
rect 544384 63106 544436 63112
rect 543004 63028 543056 63034
rect 543004 62970 543056 62976
rect 541624 62892 541676 62898
rect 541624 62834 541676 62840
rect 540336 62484 540388 62490
rect 540336 62426 540388 62432
rect 540244 62416 540296 62422
rect 540244 62358 540296 62364
rect 539600 3392 539652 3398
rect 539600 3334 539652 3340
rect 538864 2848 538916 2854
rect 538864 2790 538916 2796
rect 539612 480 539640 3334
rect 540256 2922 540284 62358
rect 540348 3194 540376 62426
rect 540796 5228 540848 5234
rect 540796 5170 540848 5176
rect 540336 3188 540388 3194
rect 540336 3130 540388 3136
rect 540244 2916 540296 2922
rect 540244 2858 540296 2864
rect 540808 480 540836 5170
rect 541636 3398 541664 62834
rect 541624 3392 541676 3398
rect 541624 3334 541676 3340
rect 543016 3330 543044 62970
rect 544292 5024 544344 5030
rect 544292 4966 544344 4972
rect 543188 3392 543240 3398
rect 543188 3334 543240 3340
rect 543004 3324 543056 3330
rect 543004 3266 543056 3272
rect 541992 2984 542044 2990
rect 541992 2926 542044 2932
rect 542004 480 542032 2926
rect 543200 480 543228 3334
rect 544304 2530 544332 4966
rect 544396 3398 544424 63106
rect 545764 62756 545816 62762
rect 545764 62698 545816 62704
rect 544384 3392 544436 3398
rect 544384 3334 544436 3340
rect 545776 3126 545804 62698
rect 546684 3324 546736 3330
rect 546684 3266 546736 3272
rect 545764 3120 545816 3126
rect 545764 3062 545816 3068
rect 545488 2848 545540 2854
rect 545488 2790 545540 2796
rect 544304 2502 544424 2530
rect 544396 480 544424 2502
rect 545500 480 545528 2790
rect 546696 480 546724 3266
rect 547156 2854 547184 63174
rect 547880 4888 547932 4894
rect 547880 4830 547932 4836
rect 547144 2848 547196 2854
rect 547144 2790 547196 2796
rect 547892 480 547920 4830
rect 548536 2990 548564 63378
rect 551284 62620 551336 62626
rect 551284 62562 551336 62568
rect 551296 3330 551324 62562
rect 555436 6866 555464 638959
rect 556816 46918 556844 639231
rect 558182 636848 558238 636857
rect 558182 636783 558238 636792
rect 556804 46912 556856 46918
rect 556804 46854 556856 46860
rect 558196 33114 558224 636783
rect 558288 525774 558316 641310
rect 562324 641028 562376 641034
rect 562324 640970 562376 640976
rect 561126 637256 561182 637265
rect 561126 637191 561182 637200
rect 560942 636984 560998 636993
rect 560942 636919 560998 636928
rect 558276 525768 558328 525774
rect 558276 525710 558328 525716
rect 558184 33108 558236 33114
rect 558184 33050 558236 33056
rect 557540 32428 557592 32434
rect 557540 32370 557592 32376
rect 557552 16574 557580 32370
rect 560956 20670 560984 636919
rect 561140 485790 561168 637191
rect 561128 485784 561180 485790
rect 561128 485726 561180 485732
rect 562336 431934 562364 640970
rect 566462 640520 566518 640529
rect 566462 640455 566518 640464
rect 565084 638240 565136 638246
rect 565084 638182 565136 638188
rect 562414 637528 562470 637537
rect 562414 637463 562470 637472
rect 562428 538218 562456 637463
rect 562416 538212 562468 538218
rect 562416 538154 562468 538160
rect 562324 431928 562376 431934
rect 562324 431870 562376 431876
rect 565096 325650 565124 638182
rect 565174 636576 565230 636585
rect 565174 636511 565230 636520
rect 565188 592006 565216 636511
rect 565176 592000 565228 592006
rect 565176 591942 565228 591948
rect 565084 325644 565136 325650
rect 565084 325586 565136 325592
rect 566476 73166 566504 640455
rect 569222 637120 569278 637129
rect 569222 637055 569278 637064
rect 569236 113150 569264 637055
rect 569328 578202 569356 641378
rect 580448 640008 580500 640014
rect 580448 639950 580500 639956
rect 580264 638852 580316 638858
rect 580264 638794 580316 638800
rect 576124 637968 576176 637974
rect 576124 637910 576176 637916
rect 574744 637832 574796 637838
rect 574744 637774 574796 637780
rect 573364 637696 573416 637702
rect 573364 637638 573416 637644
rect 569316 578196 569368 578202
rect 569316 578138 569368 578144
rect 573376 153202 573404 637638
rect 574756 193186 574784 637774
rect 576136 233238 576164 637910
rect 579712 632052 579764 632058
rect 579712 631994 579764 632000
rect 579724 630873 579752 631994
rect 579710 630864 579766 630873
rect 579710 630799 579766 630808
rect 579804 618248 579856 618254
rect 579804 618190 579856 618196
rect 579816 617545 579844 618190
rect 579802 617536 579858 617545
rect 579802 617471 579858 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 580276 258913 580304 638794
rect 580356 638716 580408 638722
rect 580356 638658 580408 638664
rect 580368 365129 580396 638658
rect 580460 418305 580488 639950
rect 580446 418296 580502 418305
rect 580446 418231 580502 418240
rect 580354 365120 580410 365129
rect 580354 365055 580410 365064
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 576124 233232 576176 233238
rect 576124 233174 576176 233180
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 574744 193180 574796 193186
rect 574744 193122 574796 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 573364 153196 573416 153202
rect 573364 153138 573416 153144
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 569224 113144 569276 113150
rect 569224 113086 569276 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 566464 73160 566516 73166
rect 566464 73102 566516 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 564532 61532 564584 61538
rect 564532 61474 564584 61480
rect 561680 61464 561732 61470
rect 561680 61406 561732 61412
rect 560944 20664 560996 20670
rect 560944 20606 560996 20612
rect 561692 16574 561720 61406
rect 564544 16574 564572 61474
rect 572812 61396 572864 61402
rect 572812 61338 572864 61344
rect 557552 16546 558592 16574
rect 561692 16546 562088 16574
rect 564544 16546 565676 16574
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 551468 4956 551520 4962
rect 551468 4898 551520 4904
rect 550272 3324 550324 3330
rect 550272 3266 550324 3272
rect 551284 3324 551336 3330
rect 551284 3266 551336 3272
rect 548524 2984 548576 2990
rect 548524 2926 548576 2932
rect 549076 2916 549128 2922
rect 549076 2858 549128 2864
rect 549088 480 549116 2858
rect 550284 480 550312 3266
rect 551480 480 551508 4898
rect 554964 4820 555016 4826
rect 554964 4762 555016 4768
rect 552664 3052 552716 3058
rect 552664 2994 552716 3000
rect 552676 480 552704 2994
rect 553768 2848 553820 2854
rect 553768 2790 553820 2796
rect 553780 480 553808 2790
rect 554976 480 555004 4762
rect 556160 4072 556212 4078
rect 556160 4014 556212 4020
rect 556172 480 556200 4014
rect 557356 2984 557408 2990
rect 557356 2926 557408 2932
rect 557368 480 557396 2926
rect 558564 480 558592 16546
rect 559748 4140 559800 4146
rect 559748 4082 559800 4088
rect 559760 480 559788 4082
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 560864 480 560892 3946
rect 562060 480 562088 16546
rect 563244 3936 563296 3942
rect 563244 3878 563296 3884
rect 563256 480 563284 3878
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 565648 480 565676 16546
rect 569132 8968 569184 8974
rect 569132 8910 569184 8916
rect 568028 3800 568080 3806
rect 568028 3742 568080 3748
rect 566832 3732 566884 3738
rect 566832 3674 566884 3680
rect 566844 480 566872 3674
rect 568040 480 568068 3742
rect 569144 480 569172 8910
rect 572824 6914 572852 61338
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 572732 6886 572852 6914
rect 571524 3664 571576 3670
rect 571524 3606 571576 3612
rect 570328 3188 570380 3194
rect 570328 3130 570380 3136
rect 570340 480 570368 3130
rect 571536 480 571564 3606
rect 572732 480 572760 6886
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 573916 3596 573968 3602
rect 573916 3538 573968 3544
rect 573928 480 573956 3538
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 577412 3392 577464 3398
rect 577412 3334 577464 3340
rect 575112 3324 575164 3330
rect 575112 3266 575164 3272
rect 575124 480 575152 3266
rect 576308 3256 576360 3262
rect 576308 3198 576360 3204
rect 576320 480 576348 3198
rect 577424 480 577452 3334
rect 578620 480 578648 3470
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582196 3120 582248 3126
rect 582196 3062 582248 3068
rect 582208 480 582236 3062
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 583404 480 583432 2994
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 4802 640736 4858 640792
rect 3422 638152 3478 638208
rect 3330 632032 3386 632088
rect 3054 606056 3110 606112
rect 3330 579944 3386 580000
rect 3330 566888 3386 566944
rect 3330 553832 3386 553888
rect 3330 527856 3386 527912
rect 3146 514800 3202 514856
rect 2962 501744 3018 501800
rect 3238 475632 3294 475688
rect 3054 462576 3110 462632
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2962 410488 3018 410544
rect 3330 397432 3386 397488
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3330 214920 3386 214976
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 2778 58520 2834 58576
rect 3606 619112 3662 619168
rect 3514 201864 3570 201920
rect 3514 188844 3516 188864
rect 3516 188844 3568 188864
rect 3568 188844 3570 188864
rect 3514 188808 3570 188844
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 11702 637608 11758 637664
rect 29642 639104 29698 639160
rect 33782 640600 33838 640656
rect 32494 636248 32550 636304
rect 33874 636384 33930 636440
rect 35254 636656 35310 636712
rect 40774 637336 40830 637392
rect 72514 640464 72570 640520
rect 68374 639240 68430 639296
rect 55862 638968 55918 639024
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 515310 640736 515366 640792
rect 511078 640600 511134 640656
rect 519450 639104 519506 639160
rect 435362 638152 435418 638208
rect 60186 637880 60242 637936
rect 64418 637880 64474 637936
rect 77022 637880 77078 637936
rect 85210 637880 85266 637936
rect 185490 637880 185546 637936
rect 198002 637880 198058 637936
rect 210514 637880 210570 637936
rect 373078 637880 373134 637936
rect 385590 637880 385646 637936
rect 398102 637880 398158 637936
rect 410614 637880 410670 637936
rect 498290 637880 498346 637936
rect 533342 637744 533398 637800
rect 556802 639240 556858 639296
rect 555422 638968 555478 639024
rect 558182 636792 558238 636848
rect 561126 637200 561182 637256
rect 560942 636928 560998 636984
rect 566462 640464 566518 640520
rect 562414 637472 562470 637528
rect 565174 636520 565230 636576
rect 569222 637064 569278 637120
rect 579710 630808 579766 630864
rect 579802 617480 579858 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 524456 580226 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 351872 580226 351928
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 579894 272176 579950 272232
rect 580446 418240 580502 418296
rect 580354 365064 580410 365120
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 4797 640794 4863 640797
rect 515305 640794 515371 640797
rect 4797 640792 515371 640794
rect 4797 640736 4802 640792
rect 4858 640736 515310 640792
rect 515366 640736 515371 640792
rect 4797 640734 515371 640736
rect 4797 640731 4863 640734
rect 515305 640731 515371 640734
rect 33777 640658 33843 640661
rect 511073 640658 511139 640661
rect 33777 640656 511139 640658
rect 33777 640600 33782 640656
rect 33838 640600 511078 640656
rect 511134 640600 511139 640656
rect 33777 640598 511139 640600
rect 33777 640595 33843 640598
rect 511073 640595 511139 640598
rect 72509 640522 72575 640525
rect 566457 640522 566523 640525
rect 72509 640520 566523 640522
rect 72509 640464 72514 640520
rect 72570 640464 566462 640520
rect 566518 640464 566523 640520
rect 72509 640462 566523 640464
rect 72509 640459 72575 640462
rect 566457 640459 566523 640462
rect 68369 639298 68435 639301
rect 556797 639298 556863 639301
rect 68369 639296 556863 639298
rect 68369 639240 68374 639296
rect 68430 639240 556802 639296
rect 556858 639240 556863 639296
rect 68369 639238 556863 639240
rect 68369 639235 68435 639238
rect 556797 639235 556863 639238
rect 29637 639162 29703 639165
rect 519445 639162 519511 639165
rect 29637 639160 519511 639162
rect 29637 639104 29642 639160
rect 29698 639104 519450 639160
rect 519506 639104 519511 639160
rect 29637 639102 519511 639104
rect 29637 639099 29703 639102
rect 519445 639099 519511 639102
rect 55857 639026 55923 639029
rect 555417 639026 555483 639029
rect 55857 639024 555483 639026
rect 55857 638968 55862 639024
rect 55918 638968 555422 639024
rect 555478 638968 555483 639024
rect 55857 638966 555483 638968
rect 55857 638963 55923 638966
rect 555417 638963 555483 638966
rect 3417 638210 3483 638213
rect 435357 638210 435423 638213
rect 3417 638208 435423 638210
rect 3417 638152 3422 638208
rect 3478 638152 435362 638208
rect 435418 638152 435423 638208
rect 3417 638150 435423 638152
rect 3417 638147 3483 638150
rect 435357 638147 435423 638150
rect 489870 638014 499590 638074
rect 60181 637940 60247 637941
rect 64413 637940 64479 637941
rect 60181 637936 60228 637940
rect 60292 637938 60298 637940
rect 60181 637880 60186 637936
rect 60181 637876 60228 637880
rect 60292 637878 60338 637938
rect 64413 637936 64460 637940
rect 64524 637938 64530 637940
rect 77017 637938 77083 637941
rect 85205 637940 85271 637941
rect 185485 637940 185551 637941
rect 197997 637940 198063 637941
rect 210509 637940 210575 637941
rect 373073 637940 373139 637941
rect 385585 637940 385651 637941
rect 398097 637940 398163 637941
rect 410609 637940 410675 637941
rect 64413 637880 64418 637936
rect 60292 637876 60298 637878
rect 64413 637876 64460 637880
rect 64524 637878 64570 637938
rect 77017 637936 84210 637938
rect 77017 637880 77022 637936
rect 77078 637880 84210 637936
rect 77017 637878 84210 637880
rect 64524 637876 64530 637878
rect 60181 637875 60247 637876
rect 64413 637875 64479 637876
rect 77017 637875 77083 637878
rect 84150 637802 84210 637878
rect 85205 637936 85252 637940
rect 85316 637938 85322 637940
rect 85205 637880 85210 637936
rect 85205 637876 85252 637880
rect 85316 637878 85362 637938
rect 185485 637936 185532 637940
rect 185596 637938 185602 637940
rect 185485 637880 185490 637936
rect 85316 637876 85322 637878
rect 185485 637876 185532 637880
rect 185596 637878 185642 637938
rect 197997 637936 198044 637940
rect 198108 637938 198114 637940
rect 197997 637880 198002 637936
rect 185596 637876 185602 637878
rect 197997 637876 198044 637880
rect 198108 637878 198154 637938
rect 210509 637936 210556 637940
rect 210620 637938 210626 637940
rect 373022 637938 373028 637940
rect 210509 637880 210514 637936
rect 198108 637876 198114 637878
rect 210509 637876 210556 637880
rect 210620 637878 210666 637938
rect 372982 637878 373028 637938
rect 373092 637936 373139 637940
rect 385534 637938 385540 637940
rect 373134 637880 373139 637936
rect 210620 637876 210626 637878
rect 373022 637876 373028 637878
rect 373092 637876 373139 637880
rect 385494 637878 385540 637938
rect 385604 637936 385651 637940
rect 398046 637938 398052 637940
rect 385646 637880 385651 637936
rect 385534 637876 385540 637878
rect 385604 637876 385651 637880
rect 398006 637878 398052 637938
rect 398116 637936 398163 637940
rect 410558 637938 410564 637940
rect 398158 637880 398163 637936
rect 398046 637876 398052 637878
rect 398116 637876 398163 637880
rect 410518 637878 410564 637938
rect 410628 637936 410675 637940
rect 410670 637880 410675 637936
rect 410558 637876 410564 637878
rect 410628 637876 410675 637880
rect 85205 637875 85271 637876
rect 185485 637875 185551 637876
rect 197997 637875 198063 637876
rect 210509 637875 210575 637876
rect 373073 637875 373139 637876
rect 385585 637875 385651 637876
rect 398097 637875 398163 637876
rect 410609 637875 410675 637876
rect 489870 637802 489930 638014
rect 498285 637938 498351 637941
rect 84150 637742 489930 637802
rect 494102 637936 498351 637938
rect 494102 637880 498290 637936
rect 498346 637880 498351 637936
rect 494102 637878 498351 637880
rect 11697 637666 11763 637669
rect 494102 637666 494162 637878
rect 498285 637875 498351 637878
rect 499530 637802 499590 638014
rect 533337 637802 533403 637805
rect 499530 637800 533403 637802
rect 499530 637744 533342 637800
rect 533398 637744 533403 637800
rect 499530 637742 533403 637744
rect 533337 637739 533403 637742
rect 11697 637664 494162 637666
rect 11697 637608 11702 637664
rect 11758 637608 494162 637664
rect 11697 637606 494162 637608
rect 11697 637603 11763 637606
rect 198038 637468 198044 637532
rect 198108 637530 198114 637532
rect 562409 637530 562475 637533
rect 198108 637470 509250 637530
rect 198108 637468 198114 637470
rect 40769 637394 40835 637397
rect 410558 637394 410564 637396
rect 40769 637392 410564 637394
rect 40769 637336 40774 637392
rect 40830 637336 410564 637392
rect 40769 637334 410564 637336
rect 40769 637331 40835 637334
rect 410558 637332 410564 637334
rect 410628 637332 410634 637396
rect 509190 637394 509250 637470
rect 528510 637528 562475 637530
rect 528510 637472 562414 637528
rect 562470 637472 562475 637528
rect 528510 637470 562475 637472
rect 528510 637394 528570 637470
rect 562409 637467 562475 637470
rect 509190 637334 528570 637394
rect 185526 637196 185532 637260
rect 185596 637258 185602 637260
rect 561121 637258 561187 637261
rect 185596 637256 561187 637258
rect 185596 637200 561126 637256
rect 561182 637200 561187 637256
rect 185596 637198 561187 637200
rect 185596 637196 185602 637198
rect 561121 637195 561187 637198
rect 85246 637060 85252 637124
rect 85316 637122 85322 637124
rect 569217 637122 569283 637125
rect 85316 637120 569283 637122
rect 85316 637064 569222 637120
rect 569278 637064 569283 637120
rect 85316 637062 569283 637064
rect 85316 637060 85322 637062
rect 569217 637059 569283 637062
rect 64454 636924 64460 636988
rect 64524 636986 64530 636988
rect 560937 636986 561003 636989
rect 64524 636984 561003 636986
rect 64524 636928 560942 636984
rect 560998 636928 561003 636984
rect 64524 636926 561003 636928
rect 64524 636924 64530 636926
rect 560937 636923 561003 636926
rect 60222 636788 60228 636852
rect 60292 636850 60298 636852
rect 558177 636850 558243 636853
rect 60292 636848 558243 636850
rect 60292 636792 558182 636848
rect 558238 636792 558243 636848
rect 60292 636790 558243 636792
rect 60292 636788 60298 636790
rect 558177 636787 558243 636790
rect 35249 636714 35315 636717
rect 398046 636714 398052 636716
rect 35249 636712 398052 636714
rect 35249 636656 35254 636712
rect 35310 636656 398052 636712
rect 35249 636654 398052 636656
rect 35249 636651 35315 636654
rect 398046 636652 398052 636654
rect 398116 636652 398122 636716
rect 210550 636516 210556 636580
rect 210620 636578 210626 636580
rect 565169 636578 565235 636581
rect 210620 636576 565235 636578
rect 210620 636520 565174 636576
rect 565230 636520 565235 636576
rect 210620 636518 565235 636520
rect 210620 636516 210626 636518
rect 565169 636515 565235 636518
rect 33869 636442 33935 636445
rect 385534 636442 385540 636444
rect 33869 636440 385540 636442
rect 33869 636384 33874 636440
rect 33930 636384 385540 636440
rect 33869 636382 385540 636384
rect 33869 636379 33935 636382
rect 385534 636380 385540 636382
rect 385604 636380 385610 636444
rect 32489 636306 32555 636309
rect 373022 636306 373028 636308
rect 32489 636304 373028 636306
rect 32489 636248 32494 636304
rect 32550 636248 373028 636304
rect 32489 636246 373028 636248
rect 32489 636243 32555 636246
rect 373022 636244 373028 636246
rect 373092 636244 373098 636308
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579705 630866 579771 630869
rect 583520 630866 584960 630956
rect 579705 630864 584960 630866
rect 579705 630808 579710 630864
rect 579766 630808 584960 630864
rect 579705 630806 584960 630808
rect 579705 630803 579771 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 579797 617538 579863 617541
rect 583520 617538 584960 617628
rect 579797 617536 584960 617538
rect 579797 617480 579802 617536
rect 579858 617480 584960 617536
rect 579797 617478 584960 617480
rect 579797 617475 579863 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3049 606114 3115 606117
rect -960 606112 3115 606114
rect -960 606056 3054 606112
rect 3110 606056 3115 606112
rect -960 606054 3115 606056
rect -960 605964 480 606054
rect 3049 606051 3115 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3141 514858 3207 514861
rect -960 514856 3207 514858
rect -960 514800 3146 514856
rect 3202 514800 3207 514856
rect -960 514798 3207 514800
rect -960 514708 480 514798
rect 3141 514795 3207 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2957 501802 3023 501805
rect -960 501800 3023 501802
rect -960 501744 2962 501800
rect 3018 501744 3023 501800
rect -960 501742 3023 501744
rect -960 501652 480 501742
rect 2957 501739 3023 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3233 475690 3299 475693
rect -960 475688 3299 475690
rect -960 475632 3238 475688
rect 3294 475632 3299 475688
rect -960 475630 3299 475632
rect -960 475540 480 475630
rect 3233 475627 3299 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580441 418298 580507 418301
rect 583520 418298 584960 418388
rect 580441 418296 584960 418298
rect 580441 418240 580446 418296
rect 580502 418240 584960 418296
rect 580441 418238 584960 418240
rect 580441 418235 580507 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580349 365122 580415 365125
rect 583520 365122 584960 365212
rect 580349 365120 584960 365122
rect 580349 365064 580354 365120
rect 580410 365064 584960 365120
rect 580349 365062 584960 365064
rect 580349 365059 580415 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2773 58578 2839 58581
rect -960 58576 2839 58578
rect -960 58520 2778 58576
rect 2834 58520 2839 58576
rect -960 58518 2839 58520
rect -960 58428 480 58518
rect 2773 58515 2839 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 60228 637936 60292 637940
rect 60228 637880 60242 637936
rect 60242 637880 60292 637936
rect 60228 637876 60292 637880
rect 64460 637936 64524 637940
rect 64460 637880 64474 637936
rect 64474 637880 64524 637936
rect 64460 637876 64524 637880
rect 85252 637936 85316 637940
rect 85252 637880 85266 637936
rect 85266 637880 85316 637936
rect 85252 637876 85316 637880
rect 185532 637936 185596 637940
rect 185532 637880 185546 637936
rect 185546 637880 185596 637936
rect 185532 637876 185596 637880
rect 198044 637936 198108 637940
rect 198044 637880 198058 637936
rect 198058 637880 198108 637936
rect 198044 637876 198108 637880
rect 210556 637936 210620 637940
rect 210556 637880 210570 637936
rect 210570 637880 210620 637936
rect 210556 637876 210620 637880
rect 373028 637936 373092 637940
rect 373028 637880 373078 637936
rect 373078 637880 373092 637936
rect 373028 637876 373092 637880
rect 385540 637936 385604 637940
rect 385540 637880 385590 637936
rect 385590 637880 385604 637936
rect 385540 637876 385604 637880
rect 398052 637936 398116 637940
rect 398052 637880 398102 637936
rect 398102 637880 398116 637936
rect 398052 637876 398116 637880
rect 410564 637936 410628 637940
rect 410564 637880 410614 637936
rect 410614 637880 410628 637936
rect 410564 637876 410628 637880
rect 198044 637468 198108 637532
rect 410564 637332 410628 637396
rect 185532 637196 185596 637260
rect 85252 637060 85316 637124
rect 64460 636924 64524 636988
rect 60228 636788 60292 636852
rect 398052 636652 398116 636716
rect 210556 636516 210620 636580
rect 385540 636380 385604 636444
rect 373028 636244 373092 636308
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 640551 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 640551 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640551 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 640551 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 640551 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 640551 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 640551 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 640551 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 640551 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 640551 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640551 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 640551 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 640551 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 640551 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 640551 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 640551 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 640551 128414 668898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 640551 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640551 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 640551 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 640551 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 640551 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 640551 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 640551 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 640551 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 640551 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640551 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 640551 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 640551 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 640551 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 640551 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 640551 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 640551 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 640551 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640551 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 640551 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 640551 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 640551 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 640551 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 640551 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 640551 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 640551 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640551 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 640551 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 640551 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 640551 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 640551 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 640551 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 640551 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 640551 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640551 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 640551 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 640551 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 640551 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 640551 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 640551 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 640551 308414 668898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 640551 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640551 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 640551 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 640551 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 640551 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 640551 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 640551 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 640551 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 640551 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640551 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 640551 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 640551 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 640551 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 640551 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 640551 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 640551 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 640551 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640551 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 640551 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 640551 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 640551 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 640551 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 640551 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 640551 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 640551 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640551 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 640551 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 640551 434414 650898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 640551 438134 654618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 640551 441854 658338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 640551 445574 662058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 640551 452414 668898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 640551 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640551 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 640551 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 640551 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 640551 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 640551 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 640551 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 640551 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 640551 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640551 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 640551 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 640551 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 640551 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 640551 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 640551 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 640551 524414 668898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 640551 528134 672618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640551 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 60227 637940 60293 637941
rect 60227 637876 60228 637940
rect 60292 637876 60293 637940
rect 60227 637875 60293 637876
rect 64459 637940 64525 637941
rect 64459 637876 64460 637940
rect 64524 637876 64525 637940
rect 64459 637875 64525 637876
rect 85251 637940 85317 637941
rect 85251 637876 85252 637940
rect 85316 637876 85317 637940
rect 85251 637875 85317 637876
rect 185531 637940 185597 637941
rect 185531 637876 185532 637940
rect 185596 637876 185597 637940
rect 185531 637875 185597 637876
rect 198043 637940 198109 637941
rect 198043 637876 198044 637940
rect 198108 637876 198109 637940
rect 198043 637875 198109 637876
rect 210555 637940 210621 637941
rect 210555 637876 210556 637940
rect 210620 637876 210621 637940
rect 210555 637875 210621 637876
rect 373027 637940 373093 637941
rect 373027 637876 373028 637940
rect 373092 637876 373093 637940
rect 373027 637875 373093 637876
rect 385539 637940 385605 637941
rect 385539 637876 385540 637940
rect 385604 637876 385605 637940
rect 385539 637875 385605 637876
rect 398051 637940 398117 637941
rect 398051 637876 398052 637940
rect 398116 637876 398117 637940
rect 398051 637875 398117 637876
rect 410563 637940 410629 637941
rect 410563 637876 410564 637940
rect 410628 637876 410629 637940
rect 410563 637875 410629 637876
rect 60230 636853 60290 637875
rect 64462 636989 64522 637875
rect 85254 637125 85314 637875
rect 185534 637261 185594 637875
rect 198046 637533 198106 637875
rect 198043 637532 198109 637533
rect 198043 637468 198044 637532
rect 198108 637468 198109 637532
rect 198043 637467 198109 637468
rect 185531 637260 185597 637261
rect 185531 637196 185532 637260
rect 185596 637196 185597 637260
rect 185531 637195 185597 637196
rect 85251 637124 85317 637125
rect 85251 637060 85252 637124
rect 85316 637060 85317 637124
rect 85251 637059 85317 637060
rect 64459 636988 64525 636989
rect 64459 636924 64460 636988
rect 64524 636924 64525 636988
rect 64459 636923 64525 636924
rect 60227 636852 60293 636853
rect 60227 636788 60228 636852
rect 60292 636788 60293 636852
rect 60227 636787 60293 636788
rect 210558 636581 210618 637875
rect 210555 636580 210621 636581
rect 210555 636516 210556 636580
rect 210620 636516 210621 636580
rect 210555 636515 210621 636516
rect 373030 636309 373090 637875
rect 385542 636445 385602 637875
rect 398054 636717 398114 637875
rect 410566 637397 410626 637875
rect 410563 637396 410629 637397
rect 410563 637332 410564 637396
rect 410628 637332 410629 637396
rect 410563 637331 410629 637332
rect 398051 636716 398117 636717
rect 398051 636652 398052 636716
rect 398116 636652 398117 636716
rect 398051 636651 398117 636652
rect 385539 636444 385605 636445
rect 385539 636380 385540 636444
rect 385604 636380 385605 636444
rect 385539 636379 385605 636380
rect 373027 636308 373093 636309
rect 373027 636244 373028 636308
rect 373092 636244 373093 636308
rect 373027 636243 373093 636244
rect 73368 633454 73688 633486
rect 73368 633218 73410 633454
rect 73646 633218 73688 633454
rect 73368 633134 73688 633218
rect 73368 632898 73410 633134
rect 73646 632898 73688 633134
rect 73368 632866 73688 632898
rect 104088 633454 104408 633486
rect 104088 633218 104130 633454
rect 104366 633218 104408 633454
rect 104088 633134 104408 633218
rect 104088 632898 104130 633134
rect 104366 632898 104408 633134
rect 104088 632866 104408 632898
rect 134808 633454 135128 633486
rect 134808 633218 134850 633454
rect 135086 633218 135128 633454
rect 134808 633134 135128 633218
rect 134808 632898 134850 633134
rect 135086 632898 135128 633134
rect 134808 632866 135128 632898
rect 165528 633454 165848 633486
rect 165528 633218 165570 633454
rect 165806 633218 165848 633454
rect 165528 633134 165848 633218
rect 165528 632898 165570 633134
rect 165806 632898 165848 633134
rect 165528 632866 165848 632898
rect 196248 633454 196568 633486
rect 196248 633218 196290 633454
rect 196526 633218 196568 633454
rect 196248 633134 196568 633218
rect 196248 632898 196290 633134
rect 196526 632898 196568 633134
rect 196248 632866 196568 632898
rect 226968 633454 227288 633486
rect 226968 633218 227010 633454
rect 227246 633218 227288 633454
rect 226968 633134 227288 633218
rect 226968 632898 227010 633134
rect 227246 632898 227288 633134
rect 226968 632866 227288 632898
rect 257688 633454 258008 633486
rect 257688 633218 257730 633454
rect 257966 633218 258008 633454
rect 257688 633134 258008 633218
rect 257688 632898 257730 633134
rect 257966 632898 258008 633134
rect 257688 632866 258008 632898
rect 288408 633454 288728 633486
rect 288408 633218 288450 633454
rect 288686 633218 288728 633454
rect 288408 633134 288728 633218
rect 288408 632898 288450 633134
rect 288686 632898 288728 633134
rect 288408 632866 288728 632898
rect 319128 633454 319448 633486
rect 319128 633218 319170 633454
rect 319406 633218 319448 633454
rect 319128 633134 319448 633218
rect 319128 632898 319170 633134
rect 319406 632898 319448 633134
rect 319128 632866 319448 632898
rect 349848 633454 350168 633486
rect 349848 633218 349890 633454
rect 350126 633218 350168 633454
rect 349848 633134 350168 633218
rect 349848 632898 349890 633134
rect 350126 632898 350168 633134
rect 349848 632866 350168 632898
rect 380568 633454 380888 633486
rect 380568 633218 380610 633454
rect 380846 633218 380888 633454
rect 380568 633134 380888 633218
rect 380568 632898 380610 633134
rect 380846 632898 380888 633134
rect 380568 632866 380888 632898
rect 411288 633454 411608 633486
rect 411288 633218 411330 633454
rect 411566 633218 411608 633454
rect 411288 633134 411608 633218
rect 411288 632898 411330 633134
rect 411566 632898 411608 633134
rect 411288 632866 411608 632898
rect 442008 633454 442328 633486
rect 442008 633218 442050 633454
rect 442286 633218 442328 633454
rect 442008 633134 442328 633218
rect 442008 632898 442050 633134
rect 442286 632898 442328 633134
rect 442008 632866 442328 632898
rect 472728 633454 473048 633486
rect 472728 633218 472770 633454
rect 473006 633218 473048 633454
rect 472728 633134 473048 633218
rect 472728 632898 472770 633134
rect 473006 632898 473048 633134
rect 472728 632866 473048 632898
rect 503448 633454 503768 633486
rect 503448 633218 503490 633454
rect 503726 633218 503768 633454
rect 503448 633134 503768 633218
rect 503448 632898 503490 633134
rect 503726 632898 503768 633134
rect 503448 632866 503768 632898
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 58008 615454 58328 615486
rect 58008 615218 58050 615454
rect 58286 615218 58328 615454
rect 58008 615134 58328 615218
rect 58008 614898 58050 615134
rect 58286 614898 58328 615134
rect 58008 614866 58328 614898
rect 88728 615454 89048 615486
rect 88728 615218 88770 615454
rect 89006 615218 89048 615454
rect 88728 615134 89048 615218
rect 88728 614898 88770 615134
rect 89006 614898 89048 615134
rect 88728 614866 89048 614898
rect 119448 615454 119768 615486
rect 119448 615218 119490 615454
rect 119726 615218 119768 615454
rect 119448 615134 119768 615218
rect 119448 614898 119490 615134
rect 119726 614898 119768 615134
rect 119448 614866 119768 614898
rect 150168 615454 150488 615486
rect 150168 615218 150210 615454
rect 150446 615218 150488 615454
rect 150168 615134 150488 615218
rect 150168 614898 150210 615134
rect 150446 614898 150488 615134
rect 150168 614866 150488 614898
rect 180888 615454 181208 615486
rect 180888 615218 180930 615454
rect 181166 615218 181208 615454
rect 180888 615134 181208 615218
rect 180888 614898 180930 615134
rect 181166 614898 181208 615134
rect 180888 614866 181208 614898
rect 211608 615454 211928 615486
rect 211608 615218 211650 615454
rect 211886 615218 211928 615454
rect 211608 615134 211928 615218
rect 211608 614898 211650 615134
rect 211886 614898 211928 615134
rect 211608 614866 211928 614898
rect 242328 615454 242648 615486
rect 242328 615218 242370 615454
rect 242606 615218 242648 615454
rect 242328 615134 242648 615218
rect 242328 614898 242370 615134
rect 242606 614898 242648 615134
rect 242328 614866 242648 614898
rect 273048 615454 273368 615486
rect 273048 615218 273090 615454
rect 273326 615218 273368 615454
rect 273048 615134 273368 615218
rect 273048 614898 273090 615134
rect 273326 614898 273368 615134
rect 273048 614866 273368 614898
rect 303768 615454 304088 615486
rect 303768 615218 303810 615454
rect 304046 615218 304088 615454
rect 303768 615134 304088 615218
rect 303768 614898 303810 615134
rect 304046 614898 304088 615134
rect 303768 614866 304088 614898
rect 334488 615454 334808 615486
rect 334488 615218 334530 615454
rect 334766 615218 334808 615454
rect 334488 615134 334808 615218
rect 334488 614898 334530 615134
rect 334766 614898 334808 615134
rect 334488 614866 334808 614898
rect 365208 615454 365528 615486
rect 365208 615218 365250 615454
rect 365486 615218 365528 615454
rect 365208 615134 365528 615218
rect 365208 614898 365250 615134
rect 365486 614898 365528 615134
rect 365208 614866 365528 614898
rect 395928 615454 396248 615486
rect 395928 615218 395970 615454
rect 396206 615218 396248 615454
rect 395928 615134 396248 615218
rect 395928 614898 395970 615134
rect 396206 614898 396248 615134
rect 395928 614866 396248 614898
rect 426648 615454 426968 615486
rect 426648 615218 426690 615454
rect 426926 615218 426968 615454
rect 426648 615134 426968 615218
rect 426648 614898 426690 615134
rect 426926 614898 426968 615134
rect 426648 614866 426968 614898
rect 457368 615454 457688 615486
rect 457368 615218 457410 615454
rect 457646 615218 457688 615454
rect 457368 615134 457688 615218
rect 457368 614898 457410 615134
rect 457646 614898 457688 615134
rect 457368 614866 457688 614898
rect 488088 615454 488408 615486
rect 488088 615218 488130 615454
rect 488366 615218 488408 615454
rect 488088 615134 488408 615218
rect 488088 614898 488130 615134
rect 488366 614898 488408 615134
rect 488088 614866 488408 614898
rect 518808 615454 519128 615486
rect 518808 615218 518850 615454
rect 519086 615218 519128 615454
rect 518808 615134 519128 615218
rect 518808 614898 518850 615134
rect 519086 614898 519128 615134
rect 518808 614866 519128 614898
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 73368 597454 73688 597486
rect 73368 597218 73410 597454
rect 73646 597218 73688 597454
rect 73368 597134 73688 597218
rect 73368 596898 73410 597134
rect 73646 596898 73688 597134
rect 73368 596866 73688 596898
rect 104088 597454 104408 597486
rect 104088 597218 104130 597454
rect 104366 597218 104408 597454
rect 104088 597134 104408 597218
rect 104088 596898 104130 597134
rect 104366 596898 104408 597134
rect 104088 596866 104408 596898
rect 134808 597454 135128 597486
rect 134808 597218 134850 597454
rect 135086 597218 135128 597454
rect 134808 597134 135128 597218
rect 134808 596898 134850 597134
rect 135086 596898 135128 597134
rect 134808 596866 135128 596898
rect 165528 597454 165848 597486
rect 165528 597218 165570 597454
rect 165806 597218 165848 597454
rect 165528 597134 165848 597218
rect 165528 596898 165570 597134
rect 165806 596898 165848 597134
rect 165528 596866 165848 596898
rect 196248 597454 196568 597486
rect 196248 597218 196290 597454
rect 196526 597218 196568 597454
rect 196248 597134 196568 597218
rect 196248 596898 196290 597134
rect 196526 596898 196568 597134
rect 196248 596866 196568 596898
rect 226968 597454 227288 597486
rect 226968 597218 227010 597454
rect 227246 597218 227288 597454
rect 226968 597134 227288 597218
rect 226968 596898 227010 597134
rect 227246 596898 227288 597134
rect 226968 596866 227288 596898
rect 257688 597454 258008 597486
rect 257688 597218 257730 597454
rect 257966 597218 258008 597454
rect 257688 597134 258008 597218
rect 257688 596898 257730 597134
rect 257966 596898 258008 597134
rect 257688 596866 258008 596898
rect 288408 597454 288728 597486
rect 288408 597218 288450 597454
rect 288686 597218 288728 597454
rect 288408 597134 288728 597218
rect 288408 596898 288450 597134
rect 288686 596898 288728 597134
rect 288408 596866 288728 596898
rect 319128 597454 319448 597486
rect 319128 597218 319170 597454
rect 319406 597218 319448 597454
rect 319128 597134 319448 597218
rect 319128 596898 319170 597134
rect 319406 596898 319448 597134
rect 319128 596866 319448 596898
rect 349848 597454 350168 597486
rect 349848 597218 349890 597454
rect 350126 597218 350168 597454
rect 349848 597134 350168 597218
rect 349848 596898 349890 597134
rect 350126 596898 350168 597134
rect 349848 596866 350168 596898
rect 380568 597454 380888 597486
rect 380568 597218 380610 597454
rect 380846 597218 380888 597454
rect 380568 597134 380888 597218
rect 380568 596898 380610 597134
rect 380846 596898 380888 597134
rect 380568 596866 380888 596898
rect 411288 597454 411608 597486
rect 411288 597218 411330 597454
rect 411566 597218 411608 597454
rect 411288 597134 411608 597218
rect 411288 596898 411330 597134
rect 411566 596898 411608 597134
rect 411288 596866 411608 596898
rect 442008 597454 442328 597486
rect 442008 597218 442050 597454
rect 442286 597218 442328 597454
rect 442008 597134 442328 597218
rect 442008 596898 442050 597134
rect 442286 596898 442328 597134
rect 442008 596866 442328 596898
rect 472728 597454 473048 597486
rect 472728 597218 472770 597454
rect 473006 597218 473048 597454
rect 472728 597134 473048 597218
rect 472728 596898 472770 597134
rect 473006 596898 473048 597134
rect 472728 596866 473048 596898
rect 503448 597454 503768 597486
rect 503448 597218 503490 597454
rect 503726 597218 503768 597454
rect 503448 597134 503768 597218
rect 503448 596898 503490 597134
rect 503726 596898 503768 597134
rect 503448 596866 503768 596898
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 58008 579454 58328 579486
rect 58008 579218 58050 579454
rect 58286 579218 58328 579454
rect 58008 579134 58328 579218
rect 58008 578898 58050 579134
rect 58286 578898 58328 579134
rect 58008 578866 58328 578898
rect 88728 579454 89048 579486
rect 88728 579218 88770 579454
rect 89006 579218 89048 579454
rect 88728 579134 89048 579218
rect 88728 578898 88770 579134
rect 89006 578898 89048 579134
rect 88728 578866 89048 578898
rect 119448 579454 119768 579486
rect 119448 579218 119490 579454
rect 119726 579218 119768 579454
rect 119448 579134 119768 579218
rect 119448 578898 119490 579134
rect 119726 578898 119768 579134
rect 119448 578866 119768 578898
rect 150168 579454 150488 579486
rect 150168 579218 150210 579454
rect 150446 579218 150488 579454
rect 150168 579134 150488 579218
rect 150168 578898 150210 579134
rect 150446 578898 150488 579134
rect 150168 578866 150488 578898
rect 180888 579454 181208 579486
rect 180888 579218 180930 579454
rect 181166 579218 181208 579454
rect 180888 579134 181208 579218
rect 180888 578898 180930 579134
rect 181166 578898 181208 579134
rect 180888 578866 181208 578898
rect 211608 579454 211928 579486
rect 211608 579218 211650 579454
rect 211886 579218 211928 579454
rect 211608 579134 211928 579218
rect 211608 578898 211650 579134
rect 211886 578898 211928 579134
rect 211608 578866 211928 578898
rect 242328 579454 242648 579486
rect 242328 579218 242370 579454
rect 242606 579218 242648 579454
rect 242328 579134 242648 579218
rect 242328 578898 242370 579134
rect 242606 578898 242648 579134
rect 242328 578866 242648 578898
rect 273048 579454 273368 579486
rect 273048 579218 273090 579454
rect 273326 579218 273368 579454
rect 273048 579134 273368 579218
rect 273048 578898 273090 579134
rect 273326 578898 273368 579134
rect 273048 578866 273368 578898
rect 303768 579454 304088 579486
rect 303768 579218 303810 579454
rect 304046 579218 304088 579454
rect 303768 579134 304088 579218
rect 303768 578898 303810 579134
rect 304046 578898 304088 579134
rect 303768 578866 304088 578898
rect 334488 579454 334808 579486
rect 334488 579218 334530 579454
rect 334766 579218 334808 579454
rect 334488 579134 334808 579218
rect 334488 578898 334530 579134
rect 334766 578898 334808 579134
rect 334488 578866 334808 578898
rect 365208 579454 365528 579486
rect 365208 579218 365250 579454
rect 365486 579218 365528 579454
rect 365208 579134 365528 579218
rect 365208 578898 365250 579134
rect 365486 578898 365528 579134
rect 365208 578866 365528 578898
rect 395928 579454 396248 579486
rect 395928 579218 395970 579454
rect 396206 579218 396248 579454
rect 395928 579134 396248 579218
rect 395928 578898 395970 579134
rect 396206 578898 396248 579134
rect 395928 578866 396248 578898
rect 426648 579454 426968 579486
rect 426648 579218 426690 579454
rect 426926 579218 426968 579454
rect 426648 579134 426968 579218
rect 426648 578898 426690 579134
rect 426926 578898 426968 579134
rect 426648 578866 426968 578898
rect 457368 579454 457688 579486
rect 457368 579218 457410 579454
rect 457646 579218 457688 579454
rect 457368 579134 457688 579218
rect 457368 578898 457410 579134
rect 457646 578898 457688 579134
rect 457368 578866 457688 578898
rect 488088 579454 488408 579486
rect 488088 579218 488130 579454
rect 488366 579218 488408 579454
rect 488088 579134 488408 579218
rect 488088 578898 488130 579134
rect 488366 578898 488408 579134
rect 488088 578866 488408 578898
rect 518808 579454 519128 579486
rect 518808 579218 518850 579454
rect 519086 579218 519128 579454
rect 518808 579134 519128 579218
rect 518808 578898 518850 579134
rect 519086 578898 519128 579134
rect 518808 578866 519128 578898
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 73368 561454 73688 561486
rect 73368 561218 73410 561454
rect 73646 561218 73688 561454
rect 73368 561134 73688 561218
rect 73368 560898 73410 561134
rect 73646 560898 73688 561134
rect 73368 560866 73688 560898
rect 104088 561454 104408 561486
rect 104088 561218 104130 561454
rect 104366 561218 104408 561454
rect 104088 561134 104408 561218
rect 104088 560898 104130 561134
rect 104366 560898 104408 561134
rect 104088 560866 104408 560898
rect 134808 561454 135128 561486
rect 134808 561218 134850 561454
rect 135086 561218 135128 561454
rect 134808 561134 135128 561218
rect 134808 560898 134850 561134
rect 135086 560898 135128 561134
rect 134808 560866 135128 560898
rect 165528 561454 165848 561486
rect 165528 561218 165570 561454
rect 165806 561218 165848 561454
rect 165528 561134 165848 561218
rect 165528 560898 165570 561134
rect 165806 560898 165848 561134
rect 165528 560866 165848 560898
rect 196248 561454 196568 561486
rect 196248 561218 196290 561454
rect 196526 561218 196568 561454
rect 196248 561134 196568 561218
rect 196248 560898 196290 561134
rect 196526 560898 196568 561134
rect 196248 560866 196568 560898
rect 226968 561454 227288 561486
rect 226968 561218 227010 561454
rect 227246 561218 227288 561454
rect 226968 561134 227288 561218
rect 226968 560898 227010 561134
rect 227246 560898 227288 561134
rect 226968 560866 227288 560898
rect 257688 561454 258008 561486
rect 257688 561218 257730 561454
rect 257966 561218 258008 561454
rect 257688 561134 258008 561218
rect 257688 560898 257730 561134
rect 257966 560898 258008 561134
rect 257688 560866 258008 560898
rect 288408 561454 288728 561486
rect 288408 561218 288450 561454
rect 288686 561218 288728 561454
rect 288408 561134 288728 561218
rect 288408 560898 288450 561134
rect 288686 560898 288728 561134
rect 288408 560866 288728 560898
rect 319128 561454 319448 561486
rect 319128 561218 319170 561454
rect 319406 561218 319448 561454
rect 319128 561134 319448 561218
rect 319128 560898 319170 561134
rect 319406 560898 319448 561134
rect 319128 560866 319448 560898
rect 349848 561454 350168 561486
rect 349848 561218 349890 561454
rect 350126 561218 350168 561454
rect 349848 561134 350168 561218
rect 349848 560898 349890 561134
rect 350126 560898 350168 561134
rect 349848 560866 350168 560898
rect 380568 561454 380888 561486
rect 380568 561218 380610 561454
rect 380846 561218 380888 561454
rect 380568 561134 380888 561218
rect 380568 560898 380610 561134
rect 380846 560898 380888 561134
rect 380568 560866 380888 560898
rect 411288 561454 411608 561486
rect 411288 561218 411330 561454
rect 411566 561218 411608 561454
rect 411288 561134 411608 561218
rect 411288 560898 411330 561134
rect 411566 560898 411608 561134
rect 411288 560866 411608 560898
rect 442008 561454 442328 561486
rect 442008 561218 442050 561454
rect 442286 561218 442328 561454
rect 442008 561134 442328 561218
rect 442008 560898 442050 561134
rect 442286 560898 442328 561134
rect 442008 560866 442328 560898
rect 472728 561454 473048 561486
rect 472728 561218 472770 561454
rect 473006 561218 473048 561454
rect 472728 561134 473048 561218
rect 472728 560898 472770 561134
rect 473006 560898 473048 561134
rect 472728 560866 473048 560898
rect 503448 561454 503768 561486
rect 503448 561218 503490 561454
rect 503726 561218 503768 561454
rect 503448 561134 503768 561218
rect 503448 560898 503490 561134
rect 503726 560898 503768 561134
rect 503448 560866 503768 560898
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 58008 543454 58328 543486
rect 58008 543218 58050 543454
rect 58286 543218 58328 543454
rect 58008 543134 58328 543218
rect 58008 542898 58050 543134
rect 58286 542898 58328 543134
rect 58008 542866 58328 542898
rect 88728 543454 89048 543486
rect 88728 543218 88770 543454
rect 89006 543218 89048 543454
rect 88728 543134 89048 543218
rect 88728 542898 88770 543134
rect 89006 542898 89048 543134
rect 88728 542866 89048 542898
rect 119448 543454 119768 543486
rect 119448 543218 119490 543454
rect 119726 543218 119768 543454
rect 119448 543134 119768 543218
rect 119448 542898 119490 543134
rect 119726 542898 119768 543134
rect 119448 542866 119768 542898
rect 150168 543454 150488 543486
rect 150168 543218 150210 543454
rect 150446 543218 150488 543454
rect 150168 543134 150488 543218
rect 150168 542898 150210 543134
rect 150446 542898 150488 543134
rect 150168 542866 150488 542898
rect 180888 543454 181208 543486
rect 180888 543218 180930 543454
rect 181166 543218 181208 543454
rect 180888 543134 181208 543218
rect 180888 542898 180930 543134
rect 181166 542898 181208 543134
rect 180888 542866 181208 542898
rect 211608 543454 211928 543486
rect 211608 543218 211650 543454
rect 211886 543218 211928 543454
rect 211608 543134 211928 543218
rect 211608 542898 211650 543134
rect 211886 542898 211928 543134
rect 211608 542866 211928 542898
rect 242328 543454 242648 543486
rect 242328 543218 242370 543454
rect 242606 543218 242648 543454
rect 242328 543134 242648 543218
rect 242328 542898 242370 543134
rect 242606 542898 242648 543134
rect 242328 542866 242648 542898
rect 273048 543454 273368 543486
rect 273048 543218 273090 543454
rect 273326 543218 273368 543454
rect 273048 543134 273368 543218
rect 273048 542898 273090 543134
rect 273326 542898 273368 543134
rect 273048 542866 273368 542898
rect 303768 543454 304088 543486
rect 303768 543218 303810 543454
rect 304046 543218 304088 543454
rect 303768 543134 304088 543218
rect 303768 542898 303810 543134
rect 304046 542898 304088 543134
rect 303768 542866 304088 542898
rect 334488 543454 334808 543486
rect 334488 543218 334530 543454
rect 334766 543218 334808 543454
rect 334488 543134 334808 543218
rect 334488 542898 334530 543134
rect 334766 542898 334808 543134
rect 334488 542866 334808 542898
rect 365208 543454 365528 543486
rect 365208 543218 365250 543454
rect 365486 543218 365528 543454
rect 365208 543134 365528 543218
rect 365208 542898 365250 543134
rect 365486 542898 365528 543134
rect 365208 542866 365528 542898
rect 395928 543454 396248 543486
rect 395928 543218 395970 543454
rect 396206 543218 396248 543454
rect 395928 543134 396248 543218
rect 395928 542898 395970 543134
rect 396206 542898 396248 543134
rect 395928 542866 396248 542898
rect 426648 543454 426968 543486
rect 426648 543218 426690 543454
rect 426926 543218 426968 543454
rect 426648 543134 426968 543218
rect 426648 542898 426690 543134
rect 426926 542898 426968 543134
rect 426648 542866 426968 542898
rect 457368 543454 457688 543486
rect 457368 543218 457410 543454
rect 457646 543218 457688 543454
rect 457368 543134 457688 543218
rect 457368 542898 457410 543134
rect 457646 542898 457688 543134
rect 457368 542866 457688 542898
rect 488088 543454 488408 543486
rect 488088 543218 488130 543454
rect 488366 543218 488408 543454
rect 488088 543134 488408 543218
rect 488088 542898 488130 543134
rect 488366 542898 488408 543134
rect 488088 542866 488408 542898
rect 518808 543454 519128 543486
rect 518808 543218 518850 543454
rect 519086 543218 519128 543454
rect 518808 543134 519128 543218
rect 518808 542898 518850 543134
rect 519086 542898 519128 543134
rect 518808 542866 519128 542898
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 73368 525454 73688 525486
rect 73368 525218 73410 525454
rect 73646 525218 73688 525454
rect 73368 525134 73688 525218
rect 73368 524898 73410 525134
rect 73646 524898 73688 525134
rect 73368 524866 73688 524898
rect 104088 525454 104408 525486
rect 104088 525218 104130 525454
rect 104366 525218 104408 525454
rect 104088 525134 104408 525218
rect 104088 524898 104130 525134
rect 104366 524898 104408 525134
rect 104088 524866 104408 524898
rect 134808 525454 135128 525486
rect 134808 525218 134850 525454
rect 135086 525218 135128 525454
rect 134808 525134 135128 525218
rect 134808 524898 134850 525134
rect 135086 524898 135128 525134
rect 134808 524866 135128 524898
rect 165528 525454 165848 525486
rect 165528 525218 165570 525454
rect 165806 525218 165848 525454
rect 165528 525134 165848 525218
rect 165528 524898 165570 525134
rect 165806 524898 165848 525134
rect 165528 524866 165848 524898
rect 196248 525454 196568 525486
rect 196248 525218 196290 525454
rect 196526 525218 196568 525454
rect 196248 525134 196568 525218
rect 196248 524898 196290 525134
rect 196526 524898 196568 525134
rect 196248 524866 196568 524898
rect 226968 525454 227288 525486
rect 226968 525218 227010 525454
rect 227246 525218 227288 525454
rect 226968 525134 227288 525218
rect 226968 524898 227010 525134
rect 227246 524898 227288 525134
rect 226968 524866 227288 524898
rect 257688 525454 258008 525486
rect 257688 525218 257730 525454
rect 257966 525218 258008 525454
rect 257688 525134 258008 525218
rect 257688 524898 257730 525134
rect 257966 524898 258008 525134
rect 257688 524866 258008 524898
rect 288408 525454 288728 525486
rect 288408 525218 288450 525454
rect 288686 525218 288728 525454
rect 288408 525134 288728 525218
rect 288408 524898 288450 525134
rect 288686 524898 288728 525134
rect 288408 524866 288728 524898
rect 319128 525454 319448 525486
rect 319128 525218 319170 525454
rect 319406 525218 319448 525454
rect 319128 525134 319448 525218
rect 319128 524898 319170 525134
rect 319406 524898 319448 525134
rect 319128 524866 319448 524898
rect 349848 525454 350168 525486
rect 349848 525218 349890 525454
rect 350126 525218 350168 525454
rect 349848 525134 350168 525218
rect 349848 524898 349890 525134
rect 350126 524898 350168 525134
rect 349848 524866 350168 524898
rect 380568 525454 380888 525486
rect 380568 525218 380610 525454
rect 380846 525218 380888 525454
rect 380568 525134 380888 525218
rect 380568 524898 380610 525134
rect 380846 524898 380888 525134
rect 380568 524866 380888 524898
rect 411288 525454 411608 525486
rect 411288 525218 411330 525454
rect 411566 525218 411608 525454
rect 411288 525134 411608 525218
rect 411288 524898 411330 525134
rect 411566 524898 411608 525134
rect 411288 524866 411608 524898
rect 442008 525454 442328 525486
rect 442008 525218 442050 525454
rect 442286 525218 442328 525454
rect 442008 525134 442328 525218
rect 442008 524898 442050 525134
rect 442286 524898 442328 525134
rect 442008 524866 442328 524898
rect 472728 525454 473048 525486
rect 472728 525218 472770 525454
rect 473006 525218 473048 525454
rect 472728 525134 473048 525218
rect 472728 524898 472770 525134
rect 473006 524898 473048 525134
rect 472728 524866 473048 524898
rect 503448 525454 503768 525486
rect 503448 525218 503490 525454
rect 503726 525218 503768 525454
rect 503448 525134 503768 525218
rect 503448 524898 503490 525134
rect 503726 524898 503768 525134
rect 503448 524866 503768 524898
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 58008 507454 58328 507486
rect 58008 507218 58050 507454
rect 58286 507218 58328 507454
rect 58008 507134 58328 507218
rect 58008 506898 58050 507134
rect 58286 506898 58328 507134
rect 58008 506866 58328 506898
rect 88728 507454 89048 507486
rect 88728 507218 88770 507454
rect 89006 507218 89048 507454
rect 88728 507134 89048 507218
rect 88728 506898 88770 507134
rect 89006 506898 89048 507134
rect 88728 506866 89048 506898
rect 119448 507454 119768 507486
rect 119448 507218 119490 507454
rect 119726 507218 119768 507454
rect 119448 507134 119768 507218
rect 119448 506898 119490 507134
rect 119726 506898 119768 507134
rect 119448 506866 119768 506898
rect 150168 507454 150488 507486
rect 150168 507218 150210 507454
rect 150446 507218 150488 507454
rect 150168 507134 150488 507218
rect 150168 506898 150210 507134
rect 150446 506898 150488 507134
rect 150168 506866 150488 506898
rect 180888 507454 181208 507486
rect 180888 507218 180930 507454
rect 181166 507218 181208 507454
rect 180888 507134 181208 507218
rect 180888 506898 180930 507134
rect 181166 506898 181208 507134
rect 180888 506866 181208 506898
rect 211608 507454 211928 507486
rect 211608 507218 211650 507454
rect 211886 507218 211928 507454
rect 211608 507134 211928 507218
rect 211608 506898 211650 507134
rect 211886 506898 211928 507134
rect 211608 506866 211928 506898
rect 242328 507454 242648 507486
rect 242328 507218 242370 507454
rect 242606 507218 242648 507454
rect 242328 507134 242648 507218
rect 242328 506898 242370 507134
rect 242606 506898 242648 507134
rect 242328 506866 242648 506898
rect 273048 507454 273368 507486
rect 273048 507218 273090 507454
rect 273326 507218 273368 507454
rect 273048 507134 273368 507218
rect 273048 506898 273090 507134
rect 273326 506898 273368 507134
rect 273048 506866 273368 506898
rect 303768 507454 304088 507486
rect 303768 507218 303810 507454
rect 304046 507218 304088 507454
rect 303768 507134 304088 507218
rect 303768 506898 303810 507134
rect 304046 506898 304088 507134
rect 303768 506866 304088 506898
rect 334488 507454 334808 507486
rect 334488 507218 334530 507454
rect 334766 507218 334808 507454
rect 334488 507134 334808 507218
rect 334488 506898 334530 507134
rect 334766 506898 334808 507134
rect 334488 506866 334808 506898
rect 365208 507454 365528 507486
rect 365208 507218 365250 507454
rect 365486 507218 365528 507454
rect 365208 507134 365528 507218
rect 365208 506898 365250 507134
rect 365486 506898 365528 507134
rect 365208 506866 365528 506898
rect 395928 507454 396248 507486
rect 395928 507218 395970 507454
rect 396206 507218 396248 507454
rect 395928 507134 396248 507218
rect 395928 506898 395970 507134
rect 396206 506898 396248 507134
rect 395928 506866 396248 506898
rect 426648 507454 426968 507486
rect 426648 507218 426690 507454
rect 426926 507218 426968 507454
rect 426648 507134 426968 507218
rect 426648 506898 426690 507134
rect 426926 506898 426968 507134
rect 426648 506866 426968 506898
rect 457368 507454 457688 507486
rect 457368 507218 457410 507454
rect 457646 507218 457688 507454
rect 457368 507134 457688 507218
rect 457368 506898 457410 507134
rect 457646 506898 457688 507134
rect 457368 506866 457688 506898
rect 488088 507454 488408 507486
rect 488088 507218 488130 507454
rect 488366 507218 488408 507454
rect 488088 507134 488408 507218
rect 488088 506898 488130 507134
rect 488366 506898 488408 507134
rect 488088 506866 488408 506898
rect 518808 507454 519128 507486
rect 518808 507218 518850 507454
rect 519086 507218 519128 507454
rect 518808 507134 519128 507218
rect 518808 506898 518850 507134
rect 519086 506898 519128 507134
rect 518808 506866 519128 506898
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 73368 489454 73688 489486
rect 73368 489218 73410 489454
rect 73646 489218 73688 489454
rect 73368 489134 73688 489218
rect 73368 488898 73410 489134
rect 73646 488898 73688 489134
rect 73368 488866 73688 488898
rect 104088 489454 104408 489486
rect 104088 489218 104130 489454
rect 104366 489218 104408 489454
rect 104088 489134 104408 489218
rect 104088 488898 104130 489134
rect 104366 488898 104408 489134
rect 104088 488866 104408 488898
rect 134808 489454 135128 489486
rect 134808 489218 134850 489454
rect 135086 489218 135128 489454
rect 134808 489134 135128 489218
rect 134808 488898 134850 489134
rect 135086 488898 135128 489134
rect 134808 488866 135128 488898
rect 165528 489454 165848 489486
rect 165528 489218 165570 489454
rect 165806 489218 165848 489454
rect 165528 489134 165848 489218
rect 165528 488898 165570 489134
rect 165806 488898 165848 489134
rect 165528 488866 165848 488898
rect 196248 489454 196568 489486
rect 196248 489218 196290 489454
rect 196526 489218 196568 489454
rect 196248 489134 196568 489218
rect 196248 488898 196290 489134
rect 196526 488898 196568 489134
rect 196248 488866 196568 488898
rect 226968 489454 227288 489486
rect 226968 489218 227010 489454
rect 227246 489218 227288 489454
rect 226968 489134 227288 489218
rect 226968 488898 227010 489134
rect 227246 488898 227288 489134
rect 226968 488866 227288 488898
rect 257688 489454 258008 489486
rect 257688 489218 257730 489454
rect 257966 489218 258008 489454
rect 257688 489134 258008 489218
rect 257688 488898 257730 489134
rect 257966 488898 258008 489134
rect 257688 488866 258008 488898
rect 288408 489454 288728 489486
rect 288408 489218 288450 489454
rect 288686 489218 288728 489454
rect 288408 489134 288728 489218
rect 288408 488898 288450 489134
rect 288686 488898 288728 489134
rect 288408 488866 288728 488898
rect 319128 489454 319448 489486
rect 319128 489218 319170 489454
rect 319406 489218 319448 489454
rect 319128 489134 319448 489218
rect 319128 488898 319170 489134
rect 319406 488898 319448 489134
rect 319128 488866 319448 488898
rect 349848 489454 350168 489486
rect 349848 489218 349890 489454
rect 350126 489218 350168 489454
rect 349848 489134 350168 489218
rect 349848 488898 349890 489134
rect 350126 488898 350168 489134
rect 349848 488866 350168 488898
rect 380568 489454 380888 489486
rect 380568 489218 380610 489454
rect 380846 489218 380888 489454
rect 380568 489134 380888 489218
rect 380568 488898 380610 489134
rect 380846 488898 380888 489134
rect 380568 488866 380888 488898
rect 411288 489454 411608 489486
rect 411288 489218 411330 489454
rect 411566 489218 411608 489454
rect 411288 489134 411608 489218
rect 411288 488898 411330 489134
rect 411566 488898 411608 489134
rect 411288 488866 411608 488898
rect 442008 489454 442328 489486
rect 442008 489218 442050 489454
rect 442286 489218 442328 489454
rect 442008 489134 442328 489218
rect 442008 488898 442050 489134
rect 442286 488898 442328 489134
rect 442008 488866 442328 488898
rect 472728 489454 473048 489486
rect 472728 489218 472770 489454
rect 473006 489218 473048 489454
rect 472728 489134 473048 489218
rect 472728 488898 472770 489134
rect 473006 488898 473048 489134
rect 472728 488866 473048 488898
rect 503448 489454 503768 489486
rect 503448 489218 503490 489454
rect 503726 489218 503768 489454
rect 503448 489134 503768 489218
rect 503448 488898 503490 489134
rect 503726 488898 503768 489134
rect 503448 488866 503768 488898
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 58008 471454 58328 471486
rect 58008 471218 58050 471454
rect 58286 471218 58328 471454
rect 58008 471134 58328 471218
rect 58008 470898 58050 471134
rect 58286 470898 58328 471134
rect 58008 470866 58328 470898
rect 88728 471454 89048 471486
rect 88728 471218 88770 471454
rect 89006 471218 89048 471454
rect 88728 471134 89048 471218
rect 88728 470898 88770 471134
rect 89006 470898 89048 471134
rect 88728 470866 89048 470898
rect 119448 471454 119768 471486
rect 119448 471218 119490 471454
rect 119726 471218 119768 471454
rect 119448 471134 119768 471218
rect 119448 470898 119490 471134
rect 119726 470898 119768 471134
rect 119448 470866 119768 470898
rect 150168 471454 150488 471486
rect 150168 471218 150210 471454
rect 150446 471218 150488 471454
rect 150168 471134 150488 471218
rect 150168 470898 150210 471134
rect 150446 470898 150488 471134
rect 150168 470866 150488 470898
rect 180888 471454 181208 471486
rect 180888 471218 180930 471454
rect 181166 471218 181208 471454
rect 180888 471134 181208 471218
rect 180888 470898 180930 471134
rect 181166 470898 181208 471134
rect 180888 470866 181208 470898
rect 211608 471454 211928 471486
rect 211608 471218 211650 471454
rect 211886 471218 211928 471454
rect 211608 471134 211928 471218
rect 211608 470898 211650 471134
rect 211886 470898 211928 471134
rect 211608 470866 211928 470898
rect 242328 471454 242648 471486
rect 242328 471218 242370 471454
rect 242606 471218 242648 471454
rect 242328 471134 242648 471218
rect 242328 470898 242370 471134
rect 242606 470898 242648 471134
rect 242328 470866 242648 470898
rect 273048 471454 273368 471486
rect 273048 471218 273090 471454
rect 273326 471218 273368 471454
rect 273048 471134 273368 471218
rect 273048 470898 273090 471134
rect 273326 470898 273368 471134
rect 273048 470866 273368 470898
rect 303768 471454 304088 471486
rect 303768 471218 303810 471454
rect 304046 471218 304088 471454
rect 303768 471134 304088 471218
rect 303768 470898 303810 471134
rect 304046 470898 304088 471134
rect 303768 470866 304088 470898
rect 334488 471454 334808 471486
rect 334488 471218 334530 471454
rect 334766 471218 334808 471454
rect 334488 471134 334808 471218
rect 334488 470898 334530 471134
rect 334766 470898 334808 471134
rect 334488 470866 334808 470898
rect 365208 471454 365528 471486
rect 365208 471218 365250 471454
rect 365486 471218 365528 471454
rect 365208 471134 365528 471218
rect 365208 470898 365250 471134
rect 365486 470898 365528 471134
rect 365208 470866 365528 470898
rect 395928 471454 396248 471486
rect 395928 471218 395970 471454
rect 396206 471218 396248 471454
rect 395928 471134 396248 471218
rect 395928 470898 395970 471134
rect 396206 470898 396248 471134
rect 395928 470866 396248 470898
rect 426648 471454 426968 471486
rect 426648 471218 426690 471454
rect 426926 471218 426968 471454
rect 426648 471134 426968 471218
rect 426648 470898 426690 471134
rect 426926 470898 426968 471134
rect 426648 470866 426968 470898
rect 457368 471454 457688 471486
rect 457368 471218 457410 471454
rect 457646 471218 457688 471454
rect 457368 471134 457688 471218
rect 457368 470898 457410 471134
rect 457646 470898 457688 471134
rect 457368 470866 457688 470898
rect 488088 471454 488408 471486
rect 488088 471218 488130 471454
rect 488366 471218 488408 471454
rect 488088 471134 488408 471218
rect 488088 470898 488130 471134
rect 488366 470898 488408 471134
rect 488088 470866 488408 470898
rect 518808 471454 519128 471486
rect 518808 471218 518850 471454
rect 519086 471218 519128 471454
rect 518808 471134 519128 471218
rect 518808 470898 518850 471134
rect 519086 470898 519128 471134
rect 518808 470866 519128 470898
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 73368 453454 73688 453486
rect 73368 453218 73410 453454
rect 73646 453218 73688 453454
rect 73368 453134 73688 453218
rect 73368 452898 73410 453134
rect 73646 452898 73688 453134
rect 73368 452866 73688 452898
rect 104088 453454 104408 453486
rect 104088 453218 104130 453454
rect 104366 453218 104408 453454
rect 104088 453134 104408 453218
rect 104088 452898 104130 453134
rect 104366 452898 104408 453134
rect 104088 452866 104408 452898
rect 134808 453454 135128 453486
rect 134808 453218 134850 453454
rect 135086 453218 135128 453454
rect 134808 453134 135128 453218
rect 134808 452898 134850 453134
rect 135086 452898 135128 453134
rect 134808 452866 135128 452898
rect 165528 453454 165848 453486
rect 165528 453218 165570 453454
rect 165806 453218 165848 453454
rect 165528 453134 165848 453218
rect 165528 452898 165570 453134
rect 165806 452898 165848 453134
rect 165528 452866 165848 452898
rect 196248 453454 196568 453486
rect 196248 453218 196290 453454
rect 196526 453218 196568 453454
rect 196248 453134 196568 453218
rect 196248 452898 196290 453134
rect 196526 452898 196568 453134
rect 196248 452866 196568 452898
rect 226968 453454 227288 453486
rect 226968 453218 227010 453454
rect 227246 453218 227288 453454
rect 226968 453134 227288 453218
rect 226968 452898 227010 453134
rect 227246 452898 227288 453134
rect 226968 452866 227288 452898
rect 257688 453454 258008 453486
rect 257688 453218 257730 453454
rect 257966 453218 258008 453454
rect 257688 453134 258008 453218
rect 257688 452898 257730 453134
rect 257966 452898 258008 453134
rect 257688 452866 258008 452898
rect 288408 453454 288728 453486
rect 288408 453218 288450 453454
rect 288686 453218 288728 453454
rect 288408 453134 288728 453218
rect 288408 452898 288450 453134
rect 288686 452898 288728 453134
rect 288408 452866 288728 452898
rect 319128 453454 319448 453486
rect 319128 453218 319170 453454
rect 319406 453218 319448 453454
rect 319128 453134 319448 453218
rect 319128 452898 319170 453134
rect 319406 452898 319448 453134
rect 319128 452866 319448 452898
rect 349848 453454 350168 453486
rect 349848 453218 349890 453454
rect 350126 453218 350168 453454
rect 349848 453134 350168 453218
rect 349848 452898 349890 453134
rect 350126 452898 350168 453134
rect 349848 452866 350168 452898
rect 380568 453454 380888 453486
rect 380568 453218 380610 453454
rect 380846 453218 380888 453454
rect 380568 453134 380888 453218
rect 380568 452898 380610 453134
rect 380846 452898 380888 453134
rect 380568 452866 380888 452898
rect 411288 453454 411608 453486
rect 411288 453218 411330 453454
rect 411566 453218 411608 453454
rect 411288 453134 411608 453218
rect 411288 452898 411330 453134
rect 411566 452898 411608 453134
rect 411288 452866 411608 452898
rect 442008 453454 442328 453486
rect 442008 453218 442050 453454
rect 442286 453218 442328 453454
rect 442008 453134 442328 453218
rect 442008 452898 442050 453134
rect 442286 452898 442328 453134
rect 442008 452866 442328 452898
rect 472728 453454 473048 453486
rect 472728 453218 472770 453454
rect 473006 453218 473048 453454
rect 472728 453134 473048 453218
rect 472728 452898 472770 453134
rect 473006 452898 473048 453134
rect 472728 452866 473048 452898
rect 503448 453454 503768 453486
rect 503448 453218 503490 453454
rect 503726 453218 503768 453454
rect 503448 453134 503768 453218
rect 503448 452898 503490 453134
rect 503726 452898 503768 453134
rect 503448 452866 503768 452898
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 58008 435454 58328 435486
rect 58008 435218 58050 435454
rect 58286 435218 58328 435454
rect 58008 435134 58328 435218
rect 58008 434898 58050 435134
rect 58286 434898 58328 435134
rect 58008 434866 58328 434898
rect 88728 435454 89048 435486
rect 88728 435218 88770 435454
rect 89006 435218 89048 435454
rect 88728 435134 89048 435218
rect 88728 434898 88770 435134
rect 89006 434898 89048 435134
rect 88728 434866 89048 434898
rect 119448 435454 119768 435486
rect 119448 435218 119490 435454
rect 119726 435218 119768 435454
rect 119448 435134 119768 435218
rect 119448 434898 119490 435134
rect 119726 434898 119768 435134
rect 119448 434866 119768 434898
rect 150168 435454 150488 435486
rect 150168 435218 150210 435454
rect 150446 435218 150488 435454
rect 150168 435134 150488 435218
rect 150168 434898 150210 435134
rect 150446 434898 150488 435134
rect 150168 434866 150488 434898
rect 180888 435454 181208 435486
rect 180888 435218 180930 435454
rect 181166 435218 181208 435454
rect 180888 435134 181208 435218
rect 180888 434898 180930 435134
rect 181166 434898 181208 435134
rect 180888 434866 181208 434898
rect 211608 435454 211928 435486
rect 211608 435218 211650 435454
rect 211886 435218 211928 435454
rect 211608 435134 211928 435218
rect 211608 434898 211650 435134
rect 211886 434898 211928 435134
rect 211608 434866 211928 434898
rect 242328 435454 242648 435486
rect 242328 435218 242370 435454
rect 242606 435218 242648 435454
rect 242328 435134 242648 435218
rect 242328 434898 242370 435134
rect 242606 434898 242648 435134
rect 242328 434866 242648 434898
rect 273048 435454 273368 435486
rect 273048 435218 273090 435454
rect 273326 435218 273368 435454
rect 273048 435134 273368 435218
rect 273048 434898 273090 435134
rect 273326 434898 273368 435134
rect 273048 434866 273368 434898
rect 303768 435454 304088 435486
rect 303768 435218 303810 435454
rect 304046 435218 304088 435454
rect 303768 435134 304088 435218
rect 303768 434898 303810 435134
rect 304046 434898 304088 435134
rect 303768 434866 304088 434898
rect 334488 435454 334808 435486
rect 334488 435218 334530 435454
rect 334766 435218 334808 435454
rect 334488 435134 334808 435218
rect 334488 434898 334530 435134
rect 334766 434898 334808 435134
rect 334488 434866 334808 434898
rect 365208 435454 365528 435486
rect 365208 435218 365250 435454
rect 365486 435218 365528 435454
rect 365208 435134 365528 435218
rect 365208 434898 365250 435134
rect 365486 434898 365528 435134
rect 365208 434866 365528 434898
rect 395928 435454 396248 435486
rect 395928 435218 395970 435454
rect 396206 435218 396248 435454
rect 395928 435134 396248 435218
rect 395928 434898 395970 435134
rect 396206 434898 396248 435134
rect 395928 434866 396248 434898
rect 426648 435454 426968 435486
rect 426648 435218 426690 435454
rect 426926 435218 426968 435454
rect 426648 435134 426968 435218
rect 426648 434898 426690 435134
rect 426926 434898 426968 435134
rect 426648 434866 426968 434898
rect 457368 435454 457688 435486
rect 457368 435218 457410 435454
rect 457646 435218 457688 435454
rect 457368 435134 457688 435218
rect 457368 434898 457410 435134
rect 457646 434898 457688 435134
rect 457368 434866 457688 434898
rect 488088 435454 488408 435486
rect 488088 435218 488130 435454
rect 488366 435218 488408 435454
rect 488088 435134 488408 435218
rect 488088 434898 488130 435134
rect 488366 434898 488408 435134
rect 488088 434866 488408 434898
rect 518808 435454 519128 435486
rect 518808 435218 518850 435454
rect 519086 435218 519128 435454
rect 518808 435134 519128 435218
rect 518808 434898 518850 435134
rect 519086 434898 519128 435134
rect 518808 434866 519128 434898
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 73368 417454 73688 417486
rect 73368 417218 73410 417454
rect 73646 417218 73688 417454
rect 73368 417134 73688 417218
rect 73368 416898 73410 417134
rect 73646 416898 73688 417134
rect 73368 416866 73688 416898
rect 104088 417454 104408 417486
rect 104088 417218 104130 417454
rect 104366 417218 104408 417454
rect 104088 417134 104408 417218
rect 104088 416898 104130 417134
rect 104366 416898 104408 417134
rect 104088 416866 104408 416898
rect 134808 417454 135128 417486
rect 134808 417218 134850 417454
rect 135086 417218 135128 417454
rect 134808 417134 135128 417218
rect 134808 416898 134850 417134
rect 135086 416898 135128 417134
rect 134808 416866 135128 416898
rect 165528 417454 165848 417486
rect 165528 417218 165570 417454
rect 165806 417218 165848 417454
rect 165528 417134 165848 417218
rect 165528 416898 165570 417134
rect 165806 416898 165848 417134
rect 165528 416866 165848 416898
rect 196248 417454 196568 417486
rect 196248 417218 196290 417454
rect 196526 417218 196568 417454
rect 196248 417134 196568 417218
rect 196248 416898 196290 417134
rect 196526 416898 196568 417134
rect 196248 416866 196568 416898
rect 226968 417454 227288 417486
rect 226968 417218 227010 417454
rect 227246 417218 227288 417454
rect 226968 417134 227288 417218
rect 226968 416898 227010 417134
rect 227246 416898 227288 417134
rect 226968 416866 227288 416898
rect 257688 417454 258008 417486
rect 257688 417218 257730 417454
rect 257966 417218 258008 417454
rect 257688 417134 258008 417218
rect 257688 416898 257730 417134
rect 257966 416898 258008 417134
rect 257688 416866 258008 416898
rect 288408 417454 288728 417486
rect 288408 417218 288450 417454
rect 288686 417218 288728 417454
rect 288408 417134 288728 417218
rect 288408 416898 288450 417134
rect 288686 416898 288728 417134
rect 288408 416866 288728 416898
rect 319128 417454 319448 417486
rect 319128 417218 319170 417454
rect 319406 417218 319448 417454
rect 319128 417134 319448 417218
rect 319128 416898 319170 417134
rect 319406 416898 319448 417134
rect 319128 416866 319448 416898
rect 349848 417454 350168 417486
rect 349848 417218 349890 417454
rect 350126 417218 350168 417454
rect 349848 417134 350168 417218
rect 349848 416898 349890 417134
rect 350126 416898 350168 417134
rect 349848 416866 350168 416898
rect 380568 417454 380888 417486
rect 380568 417218 380610 417454
rect 380846 417218 380888 417454
rect 380568 417134 380888 417218
rect 380568 416898 380610 417134
rect 380846 416898 380888 417134
rect 380568 416866 380888 416898
rect 411288 417454 411608 417486
rect 411288 417218 411330 417454
rect 411566 417218 411608 417454
rect 411288 417134 411608 417218
rect 411288 416898 411330 417134
rect 411566 416898 411608 417134
rect 411288 416866 411608 416898
rect 442008 417454 442328 417486
rect 442008 417218 442050 417454
rect 442286 417218 442328 417454
rect 442008 417134 442328 417218
rect 442008 416898 442050 417134
rect 442286 416898 442328 417134
rect 442008 416866 442328 416898
rect 472728 417454 473048 417486
rect 472728 417218 472770 417454
rect 473006 417218 473048 417454
rect 472728 417134 473048 417218
rect 472728 416898 472770 417134
rect 473006 416898 473048 417134
rect 472728 416866 473048 416898
rect 503448 417454 503768 417486
rect 503448 417218 503490 417454
rect 503726 417218 503768 417454
rect 503448 417134 503768 417218
rect 503448 416898 503490 417134
rect 503726 416898 503768 417134
rect 503448 416866 503768 416898
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 58008 399454 58328 399486
rect 58008 399218 58050 399454
rect 58286 399218 58328 399454
rect 58008 399134 58328 399218
rect 58008 398898 58050 399134
rect 58286 398898 58328 399134
rect 58008 398866 58328 398898
rect 88728 399454 89048 399486
rect 88728 399218 88770 399454
rect 89006 399218 89048 399454
rect 88728 399134 89048 399218
rect 88728 398898 88770 399134
rect 89006 398898 89048 399134
rect 88728 398866 89048 398898
rect 119448 399454 119768 399486
rect 119448 399218 119490 399454
rect 119726 399218 119768 399454
rect 119448 399134 119768 399218
rect 119448 398898 119490 399134
rect 119726 398898 119768 399134
rect 119448 398866 119768 398898
rect 150168 399454 150488 399486
rect 150168 399218 150210 399454
rect 150446 399218 150488 399454
rect 150168 399134 150488 399218
rect 150168 398898 150210 399134
rect 150446 398898 150488 399134
rect 150168 398866 150488 398898
rect 180888 399454 181208 399486
rect 180888 399218 180930 399454
rect 181166 399218 181208 399454
rect 180888 399134 181208 399218
rect 180888 398898 180930 399134
rect 181166 398898 181208 399134
rect 180888 398866 181208 398898
rect 211608 399454 211928 399486
rect 211608 399218 211650 399454
rect 211886 399218 211928 399454
rect 211608 399134 211928 399218
rect 211608 398898 211650 399134
rect 211886 398898 211928 399134
rect 211608 398866 211928 398898
rect 242328 399454 242648 399486
rect 242328 399218 242370 399454
rect 242606 399218 242648 399454
rect 242328 399134 242648 399218
rect 242328 398898 242370 399134
rect 242606 398898 242648 399134
rect 242328 398866 242648 398898
rect 273048 399454 273368 399486
rect 273048 399218 273090 399454
rect 273326 399218 273368 399454
rect 273048 399134 273368 399218
rect 273048 398898 273090 399134
rect 273326 398898 273368 399134
rect 273048 398866 273368 398898
rect 303768 399454 304088 399486
rect 303768 399218 303810 399454
rect 304046 399218 304088 399454
rect 303768 399134 304088 399218
rect 303768 398898 303810 399134
rect 304046 398898 304088 399134
rect 303768 398866 304088 398898
rect 334488 399454 334808 399486
rect 334488 399218 334530 399454
rect 334766 399218 334808 399454
rect 334488 399134 334808 399218
rect 334488 398898 334530 399134
rect 334766 398898 334808 399134
rect 334488 398866 334808 398898
rect 365208 399454 365528 399486
rect 365208 399218 365250 399454
rect 365486 399218 365528 399454
rect 365208 399134 365528 399218
rect 365208 398898 365250 399134
rect 365486 398898 365528 399134
rect 365208 398866 365528 398898
rect 395928 399454 396248 399486
rect 395928 399218 395970 399454
rect 396206 399218 396248 399454
rect 395928 399134 396248 399218
rect 395928 398898 395970 399134
rect 396206 398898 396248 399134
rect 395928 398866 396248 398898
rect 426648 399454 426968 399486
rect 426648 399218 426690 399454
rect 426926 399218 426968 399454
rect 426648 399134 426968 399218
rect 426648 398898 426690 399134
rect 426926 398898 426968 399134
rect 426648 398866 426968 398898
rect 457368 399454 457688 399486
rect 457368 399218 457410 399454
rect 457646 399218 457688 399454
rect 457368 399134 457688 399218
rect 457368 398898 457410 399134
rect 457646 398898 457688 399134
rect 457368 398866 457688 398898
rect 488088 399454 488408 399486
rect 488088 399218 488130 399454
rect 488366 399218 488408 399454
rect 488088 399134 488408 399218
rect 488088 398898 488130 399134
rect 488366 398898 488408 399134
rect 488088 398866 488408 398898
rect 518808 399454 519128 399486
rect 518808 399218 518850 399454
rect 519086 399218 519128 399454
rect 518808 399134 519128 399218
rect 518808 398898 518850 399134
rect 519086 398898 519128 399134
rect 518808 398866 519128 398898
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 73368 381454 73688 381486
rect 73368 381218 73410 381454
rect 73646 381218 73688 381454
rect 73368 381134 73688 381218
rect 73368 380898 73410 381134
rect 73646 380898 73688 381134
rect 73368 380866 73688 380898
rect 104088 381454 104408 381486
rect 104088 381218 104130 381454
rect 104366 381218 104408 381454
rect 104088 381134 104408 381218
rect 104088 380898 104130 381134
rect 104366 380898 104408 381134
rect 104088 380866 104408 380898
rect 134808 381454 135128 381486
rect 134808 381218 134850 381454
rect 135086 381218 135128 381454
rect 134808 381134 135128 381218
rect 134808 380898 134850 381134
rect 135086 380898 135128 381134
rect 134808 380866 135128 380898
rect 165528 381454 165848 381486
rect 165528 381218 165570 381454
rect 165806 381218 165848 381454
rect 165528 381134 165848 381218
rect 165528 380898 165570 381134
rect 165806 380898 165848 381134
rect 165528 380866 165848 380898
rect 196248 381454 196568 381486
rect 196248 381218 196290 381454
rect 196526 381218 196568 381454
rect 196248 381134 196568 381218
rect 196248 380898 196290 381134
rect 196526 380898 196568 381134
rect 196248 380866 196568 380898
rect 226968 381454 227288 381486
rect 226968 381218 227010 381454
rect 227246 381218 227288 381454
rect 226968 381134 227288 381218
rect 226968 380898 227010 381134
rect 227246 380898 227288 381134
rect 226968 380866 227288 380898
rect 257688 381454 258008 381486
rect 257688 381218 257730 381454
rect 257966 381218 258008 381454
rect 257688 381134 258008 381218
rect 257688 380898 257730 381134
rect 257966 380898 258008 381134
rect 257688 380866 258008 380898
rect 288408 381454 288728 381486
rect 288408 381218 288450 381454
rect 288686 381218 288728 381454
rect 288408 381134 288728 381218
rect 288408 380898 288450 381134
rect 288686 380898 288728 381134
rect 288408 380866 288728 380898
rect 319128 381454 319448 381486
rect 319128 381218 319170 381454
rect 319406 381218 319448 381454
rect 319128 381134 319448 381218
rect 319128 380898 319170 381134
rect 319406 380898 319448 381134
rect 319128 380866 319448 380898
rect 349848 381454 350168 381486
rect 349848 381218 349890 381454
rect 350126 381218 350168 381454
rect 349848 381134 350168 381218
rect 349848 380898 349890 381134
rect 350126 380898 350168 381134
rect 349848 380866 350168 380898
rect 380568 381454 380888 381486
rect 380568 381218 380610 381454
rect 380846 381218 380888 381454
rect 380568 381134 380888 381218
rect 380568 380898 380610 381134
rect 380846 380898 380888 381134
rect 380568 380866 380888 380898
rect 411288 381454 411608 381486
rect 411288 381218 411330 381454
rect 411566 381218 411608 381454
rect 411288 381134 411608 381218
rect 411288 380898 411330 381134
rect 411566 380898 411608 381134
rect 411288 380866 411608 380898
rect 442008 381454 442328 381486
rect 442008 381218 442050 381454
rect 442286 381218 442328 381454
rect 442008 381134 442328 381218
rect 442008 380898 442050 381134
rect 442286 380898 442328 381134
rect 442008 380866 442328 380898
rect 472728 381454 473048 381486
rect 472728 381218 472770 381454
rect 473006 381218 473048 381454
rect 472728 381134 473048 381218
rect 472728 380898 472770 381134
rect 473006 380898 473048 381134
rect 472728 380866 473048 380898
rect 503448 381454 503768 381486
rect 503448 381218 503490 381454
rect 503726 381218 503768 381454
rect 503448 381134 503768 381218
rect 503448 380898 503490 381134
rect 503726 380898 503768 381134
rect 503448 380866 503768 380898
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 58008 363454 58328 363486
rect 58008 363218 58050 363454
rect 58286 363218 58328 363454
rect 58008 363134 58328 363218
rect 58008 362898 58050 363134
rect 58286 362898 58328 363134
rect 58008 362866 58328 362898
rect 88728 363454 89048 363486
rect 88728 363218 88770 363454
rect 89006 363218 89048 363454
rect 88728 363134 89048 363218
rect 88728 362898 88770 363134
rect 89006 362898 89048 363134
rect 88728 362866 89048 362898
rect 119448 363454 119768 363486
rect 119448 363218 119490 363454
rect 119726 363218 119768 363454
rect 119448 363134 119768 363218
rect 119448 362898 119490 363134
rect 119726 362898 119768 363134
rect 119448 362866 119768 362898
rect 150168 363454 150488 363486
rect 150168 363218 150210 363454
rect 150446 363218 150488 363454
rect 150168 363134 150488 363218
rect 150168 362898 150210 363134
rect 150446 362898 150488 363134
rect 150168 362866 150488 362898
rect 180888 363454 181208 363486
rect 180888 363218 180930 363454
rect 181166 363218 181208 363454
rect 180888 363134 181208 363218
rect 180888 362898 180930 363134
rect 181166 362898 181208 363134
rect 180888 362866 181208 362898
rect 211608 363454 211928 363486
rect 211608 363218 211650 363454
rect 211886 363218 211928 363454
rect 211608 363134 211928 363218
rect 211608 362898 211650 363134
rect 211886 362898 211928 363134
rect 211608 362866 211928 362898
rect 242328 363454 242648 363486
rect 242328 363218 242370 363454
rect 242606 363218 242648 363454
rect 242328 363134 242648 363218
rect 242328 362898 242370 363134
rect 242606 362898 242648 363134
rect 242328 362866 242648 362898
rect 273048 363454 273368 363486
rect 273048 363218 273090 363454
rect 273326 363218 273368 363454
rect 273048 363134 273368 363218
rect 273048 362898 273090 363134
rect 273326 362898 273368 363134
rect 273048 362866 273368 362898
rect 303768 363454 304088 363486
rect 303768 363218 303810 363454
rect 304046 363218 304088 363454
rect 303768 363134 304088 363218
rect 303768 362898 303810 363134
rect 304046 362898 304088 363134
rect 303768 362866 304088 362898
rect 334488 363454 334808 363486
rect 334488 363218 334530 363454
rect 334766 363218 334808 363454
rect 334488 363134 334808 363218
rect 334488 362898 334530 363134
rect 334766 362898 334808 363134
rect 334488 362866 334808 362898
rect 365208 363454 365528 363486
rect 365208 363218 365250 363454
rect 365486 363218 365528 363454
rect 365208 363134 365528 363218
rect 365208 362898 365250 363134
rect 365486 362898 365528 363134
rect 365208 362866 365528 362898
rect 395928 363454 396248 363486
rect 395928 363218 395970 363454
rect 396206 363218 396248 363454
rect 395928 363134 396248 363218
rect 395928 362898 395970 363134
rect 396206 362898 396248 363134
rect 395928 362866 396248 362898
rect 426648 363454 426968 363486
rect 426648 363218 426690 363454
rect 426926 363218 426968 363454
rect 426648 363134 426968 363218
rect 426648 362898 426690 363134
rect 426926 362898 426968 363134
rect 426648 362866 426968 362898
rect 457368 363454 457688 363486
rect 457368 363218 457410 363454
rect 457646 363218 457688 363454
rect 457368 363134 457688 363218
rect 457368 362898 457410 363134
rect 457646 362898 457688 363134
rect 457368 362866 457688 362898
rect 488088 363454 488408 363486
rect 488088 363218 488130 363454
rect 488366 363218 488408 363454
rect 488088 363134 488408 363218
rect 488088 362898 488130 363134
rect 488366 362898 488408 363134
rect 488088 362866 488408 362898
rect 518808 363454 519128 363486
rect 518808 363218 518850 363454
rect 519086 363218 519128 363454
rect 518808 363134 519128 363218
rect 518808 362898 518850 363134
rect 519086 362898 519128 363134
rect 518808 362866 519128 362898
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 73368 345454 73688 345486
rect 73368 345218 73410 345454
rect 73646 345218 73688 345454
rect 73368 345134 73688 345218
rect 73368 344898 73410 345134
rect 73646 344898 73688 345134
rect 73368 344866 73688 344898
rect 104088 345454 104408 345486
rect 104088 345218 104130 345454
rect 104366 345218 104408 345454
rect 104088 345134 104408 345218
rect 104088 344898 104130 345134
rect 104366 344898 104408 345134
rect 104088 344866 104408 344898
rect 134808 345454 135128 345486
rect 134808 345218 134850 345454
rect 135086 345218 135128 345454
rect 134808 345134 135128 345218
rect 134808 344898 134850 345134
rect 135086 344898 135128 345134
rect 134808 344866 135128 344898
rect 165528 345454 165848 345486
rect 165528 345218 165570 345454
rect 165806 345218 165848 345454
rect 165528 345134 165848 345218
rect 165528 344898 165570 345134
rect 165806 344898 165848 345134
rect 165528 344866 165848 344898
rect 196248 345454 196568 345486
rect 196248 345218 196290 345454
rect 196526 345218 196568 345454
rect 196248 345134 196568 345218
rect 196248 344898 196290 345134
rect 196526 344898 196568 345134
rect 196248 344866 196568 344898
rect 226968 345454 227288 345486
rect 226968 345218 227010 345454
rect 227246 345218 227288 345454
rect 226968 345134 227288 345218
rect 226968 344898 227010 345134
rect 227246 344898 227288 345134
rect 226968 344866 227288 344898
rect 257688 345454 258008 345486
rect 257688 345218 257730 345454
rect 257966 345218 258008 345454
rect 257688 345134 258008 345218
rect 257688 344898 257730 345134
rect 257966 344898 258008 345134
rect 257688 344866 258008 344898
rect 288408 345454 288728 345486
rect 288408 345218 288450 345454
rect 288686 345218 288728 345454
rect 288408 345134 288728 345218
rect 288408 344898 288450 345134
rect 288686 344898 288728 345134
rect 288408 344866 288728 344898
rect 319128 345454 319448 345486
rect 319128 345218 319170 345454
rect 319406 345218 319448 345454
rect 319128 345134 319448 345218
rect 319128 344898 319170 345134
rect 319406 344898 319448 345134
rect 319128 344866 319448 344898
rect 349848 345454 350168 345486
rect 349848 345218 349890 345454
rect 350126 345218 350168 345454
rect 349848 345134 350168 345218
rect 349848 344898 349890 345134
rect 350126 344898 350168 345134
rect 349848 344866 350168 344898
rect 380568 345454 380888 345486
rect 380568 345218 380610 345454
rect 380846 345218 380888 345454
rect 380568 345134 380888 345218
rect 380568 344898 380610 345134
rect 380846 344898 380888 345134
rect 380568 344866 380888 344898
rect 411288 345454 411608 345486
rect 411288 345218 411330 345454
rect 411566 345218 411608 345454
rect 411288 345134 411608 345218
rect 411288 344898 411330 345134
rect 411566 344898 411608 345134
rect 411288 344866 411608 344898
rect 442008 345454 442328 345486
rect 442008 345218 442050 345454
rect 442286 345218 442328 345454
rect 442008 345134 442328 345218
rect 442008 344898 442050 345134
rect 442286 344898 442328 345134
rect 442008 344866 442328 344898
rect 472728 345454 473048 345486
rect 472728 345218 472770 345454
rect 473006 345218 473048 345454
rect 472728 345134 473048 345218
rect 472728 344898 472770 345134
rect 473006 344898 473048 345134
rect 472728 344866 473048 344898
rect 503448 345454 503768 345486
rect 503448 345218 503490 345454
rect 503726 345218 503768 345454
rect 503448 345134 503768 345218
rect 503448 344898 503490 345134
rect 503726 344898 503768 345134
rect 503448 344866 503768 344898
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 58008 327454 58328 327486
rect 58008 327218 58050 327454
rect 58286 327218 58328 327454
rect 58008 327134 58328 327218
rect 58008 326898 58050 327134
rect 58286 326898 58328 327134
rect 58008 326866 58328 326898
rect 88728 327454 89048 327486
rect 88728 327218 88770 327454
rect 89006 327218 89048 327454
rect 88728 327134 89048 327218
rect 88728 326898 88770 327134
rect 89006 326898 89048 327134
rect 88728 326866 89048 326898
rect 119448 327454 119768 327486
rect 119448 327218 119490 327454
rect 119726 327218 119768 327454
rect 119448 327134 119768 327218
rect 119448 326898 119490 327134
rect 119726 326898 119768 327134
rect 119448 326866 119768 326898
rect 150168 327454 150488 327486
rect 150168 327218 150210 327454
rect 150446 327218 150488 327454
rect 150168 327134 150488 327218
rect 150168 326898 150210 327134
rect 150446 326898 150488 327134
rect 150168 326866 150488 326898
rect 180888 327454 181208 327486
rect 180888 327218 180930 327454
rect 181166 327218 181208 327454
rect 180888 327134 181208 327218
rect 180888 326898 180930 327134
rect 181166 326898 181208 327134
rect 180888 326866 181208 326898
rect 211608 327454 211928 327486
rect 211608 327218 211650 327454
rect 211886 327218 211928 327454
rect 211608 327134 211928 327218
rect 211608 326898 211650 327134
rect 211886 326898 211928 327134
rect 211608 326866 211928 326898
rect 242328 327454 242648 327486
rect 242328 327218 242370 327454
rect 242606 327218 242648 327454
rect 242328 327134 242648 327218
rect 242328 326898 242370 327134
rect 242606 326898 242648 327134
rect 242328 326866 242648 326898
rect 273048 327454 273368 327486
rect 273048 327218 273090 327454
rect 273326 327218 273368 327454
rect 273048 327134 273368 327218
rect 273048 326898 273090 327134
rect 273326 326898 273368 327134
rect 273048 326866 273368 326898
rect 303768 327454 304088 327486
rect 303768 327218 303810 327454
rect 304046 327218 304088 327454
rect 303768 327134 304088 327218
rect 303768 326898 303810 327134
rect 304046 326898 304088 327134
rect 303768 326866 304088 326898
rect 334488 327454 334808 327486
rect 334488 327218 334530 327454
rect 334766 327218 334808 327454
rect 334488 327134 334808 327218
rect 334488 326898 334530 327134
rect 334766 326898 334808 327134
rect 334488 326866 334808 326898
rect 365208 327454 365528 327486
rect 365208 327218 365250 327454
rect 365486 327218 365528 327454
rect 365208 327134 365528 327218
rect 365208 326898 365250 327134
rect 365486 326898 365528 327134
rect 365208 326866 365528 326898
rect 395928 327454 396248 327486
rect 395928 327218 395970 327454
rect 396206 327218 396248 327454
rect 395928 327134 396248 327218
rect 395928 326898 395970 327134
rect 396206 326898 396248 327134
rect 395928 326866 396248 326898
rect 426648 327454 426968 327486
rect 426648 327218 426690 327454
rect 426926 327218 426968 327454
rect 426648 327134 426968 327218
rect 426648 326898 426690 327134
rect 426926 326898 426968 327134
rect 426648 326866 426968 326898
rect 457368 327454 457688 327486
rect 457368 327218 457410 327454
rect 457646 327218 457688 327454
rect 457368 327134 457688 327218
rect 457368 326898 457410 327134
rect 457646 326898 457688 327134
rect 457368 326866 457688 326898
rect 488088 327454 488408 327486
rect 488088 327218 488130 327454
rect 488366 327218 488408 327454
rect 488088 327134 488408 327218
rect 488088 326898 488130 327134
rect 488366 326898 488408 327134
rect 488088 326866 488408 326898
rect 518808 327454 519128 327486
rect 518808 327218 518850 327454
rect 519086 327218 519128 327454
rect 518808 327134 519128 327218
rect 518808 326898 518850 327134
rect 519086 326898 519128 327134
rect 518808 326866 519128 326898
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 73368 309454 73688 309486
rect 73368 309218 73410 309454
rect 73646 309218 73688 309454
rect 73368 309134 73688 309218
rect 73368 308898 73410 309134
rect 73646 308898 73688 309134
rect 73368 308866 73688 308898
rect 104088 309454 104408 309486
rect 104088 309218 104130 309454
rect 104366 309218 104408 309454
rect 104088 309134 104408 309218
rect 104088 308898 104130 309134
rect 104366 308898 104408 309134
rect 104088 308866 104408 308898
rect 134808 309454 135128 309486
rect 134808 309218 134850 309454
rect 135086 309218 135128 309454
rect 134808 309134 135128 309218
rect 134808 308898 134850 309134
rect 135086 308898 135128 309134
rect 134808 308866 135128 308898
rect 165528 309454 165848 309486
rect 165528 309218 165570 309454
rect 165806 309218 165848 309454
rect 165528 309134 165848 309218
rect 165528 308898 165570 309134
rect 165806 308898 165848 309134
rect 165528 308866 165848 308898
rect 196248 309454 196568 309486
rect 196248 309218 196290 309454
rect 196526 309218 196568 309454
rect 196248 309134 196568 309218
rect 196248 308898 196290 309134
rect 196526 308898 196568 309134
rect 196248 308866 196568 308898
rect 226968 309454 227288 309486
rect 226968 309218 227010 309454
rect 227246 309218 227288 309454
rect 226968 309134 227288 309218
rect 226968 308898 227010 309134
rect 227246 308898 227288 309134
rect 226968 308866 227288 308898
rect 257688 309454 258008 309486
rect 257688 309218 257730 309454
rect 257966 309218 258008 309454
rect 257688 309134 258008 309218
rect 257688 308898 257730 309134
rect 257966 308898 258008 309134
rect 257688 308866 258008 308898
rect 288408 309454 288728 309486
rect 288408 309218 288450 309454
rect 288686 309218 288728 309454
rect 288408 309134 288728 309218
rect 288408 308898 288450 309134
rect 288686 308898 288728 309134
rect 288408 308866 288728 308898
rect 319128 309454 319448 309486
rect 319128 309218 319170 309454
rect 319406 309218 319448 309454
rect 319128 309134 319448 309218
rect 319128 308898 319170 309134
rect 319406 308898 319448 309134
rect 319128 308866 319448 308898
rect 349848 309454 350168 309486
rect 349848 309218 349890 309454
rect 350126 309218 350168 309454
rect 349848 309134 350168 309218
rect 349848 308898 349890 309134
rect 350126 308898 350168 309134
rect 349848 308866 350168 308898
rect 380568 309454 380888 309486
rect 380568 309218 380610 309454
rect 380846 309218 380888 309454
rect 380568 309134 380888 309218
rect 380568 308898 380610 309134
rect 380846 308898 380888 309134
rect 380568 308866 380888 308898
rect 411288 309454 411608 309486
rect 411288 309218 411330 309454
rect 411566 309218 411608 309454
rect 411288 309134 411608 309218
rect 411288 308898 411330 309134
rect 411566 308898 411608 309134
rect 411288 308866 411608 308898
rect 442008 309454 442328 309486
rect 442008 309218 442050 309454
rect 442286 309218 442328 309454
rect 442008 309134 442328 309218
rect 442008 308898 442050 309134
rect 442286 308898 442328 309134
rect 442008 308866 442328 308898
rect 472728 309454 473048 309486
rect 472728 309218 472770 309454
rect 473006 309218 473048 309454
rect 472728 309134 473048 309218
rect 472728 308898 472770 309134
rect 473006 308898 473048 309134
rect 472728 308866 473048 308898
rect 503448 309454 503768 309486
rect 503448 309218 503490 309454
rect 503726 309218 503768 309454
rect 503448 309134 503768 309218
rect 503448 308898 503490 309134
rect 503726 308898 503768 309134
rect 503448 308866 503768 308898
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 58008 291454 58328 291486
rect 58008 291218 58050 291454
rect 58286 291218 58328 291454
rect 58008 291134 58328 291218
rect 58008 290898 58050 291134
rect 58286 290898 58328 291134
rect 58008 290866 58328 290898
rect 88728 291454 89048 291486
rect 88728 291218 88770 291454
rect 89006 291218 89048 291454
rect 88728 291134 89048 291218
rect 88728 290898 88770 291134
rect 89006 290898 89048 291134
rect 88728 290866 89048 290898
rect 119448 291454 119768 291486
rect 119448 291218 119490 291454
rect 119726 291218 119768 291454
rect 119448 291134 119768 291218
rect 119448 290898 119490 291134
rect 119726 290898 119768 291134
rect 119448 290866 119768 290898
rect 150168 291454 150488 291486
rect 150168 291218 150210 291454
rect 150446 291218 150488 291454
rect 150168 291134 150488 291218
rect 150168 290898 150210 291134
rect 150446 290898 150488 291134
rect 150168 290866 150488 290898
rect 180888 291454 181208 291486
rect 180888 291218 180930 291454
rect 181166 291218 181208 291454
rect 180888 291134 181208 291218
rect 180888 290898 180930 291134
rect 181166 290898 181208 291134
rect 180888 290866 181208 290898
rect 211608 291454 211928 291486
rect 211608 291218 211650 291454
rect 211886 291218 211928 291454
rect 211608 291134 211928 291218
rect 211608 290898 211650 291134
rect 211886 290898 211928 291134
rect 211608 290866 211928 290898
rect 242328 291454 242648 291486
rect 242328 291218 242370 291454
rect 242606 291218 242648 291454
rect 242328 291134 242648 291218
rect 242328 290898 242370 291134
rect 242606 290898 242648 291134
rect 242328 290866 242648 290898
rect 273048 291454 273368 291486
rect 273048 291218 273090 291454
rect 273326 291218 273368 291454
rect 273048 291134 273368 291218
rect 273048 290898 273090 291134
rect 273326 290898 273368 291134
rect 273048 290866 273368 290898
rect 303768 291454 304088 291486
rect 303768 291218 303810 291454
rect 304046 291218 304088 291454
rect 303768 291134 304088 291218
rect 303768 290898 303810 291134
rect 304046 290898 304088 291134
rect 303768 290866 304088 290898
rect 334488 291454 334808 291486
rect 334488 291218 334530 291454
rect 334766 291218 334808 291454
rect 334488 291134 334808 291218
rect 334488 290898 334530 291134
rect 334766 290898 334808 291134
rect 334488 290866 334808 290898
rect 365208 291454 365528 291486
rect 365208 291218 365250 291454
rect 365486 291218 365528 291454
rect 365208 291134 365528 291218
rect 365208 290898 365250 291134
rect 365486 290898 365528 291134
rect 365208 290866 365528 290898
rect 395928 291454 396248 291486
rect 395928 291218 395970 291454
rect 396206 291218 396248 291454
rect 395928 291134 396248 291218
rect 395928 290898 395970 291134
rect 396206 290898 396248 291134
rect 395928 290866 396248 290898
rect 426648 291454 426968 291486
rect 426648 291218 426690 291454
rect 426926 291218 426968 291454
rect 426648 291134 426968 291218
rect 426648 290898 426690 291134
rect 426926 290898 426968 291134
rect 426648 290866 426968 290898
rect 457368 291454 457688 291486
rect 457368 291218 457410 291454
rect 457646 291218 457688 291454
rect 457368 291134 457688 291218
rect 457368 290898 457410 291134
rect 457646 290898 457688 291134
rect 457368 290866 457688 290898
rect 488088 291454 488408 291486
rect 488088 291218 488130 291454
rect 488366 291218 488408 291454
rect 488088 291134 488408 291218
rect 488088 290898 488130 291134
rect 488366 290898 488408 291134
rect 488088 290866 488408 290898
rect 518808 291454 519128 291486
rect 518808 291218 518850 291454
rect 519086 291218 519128 291454
rect 518808 291134 519128 291218
rect 518808 290898 518850 291134
rect 519086 290898 519128 291134
rect 518808 290866 519128 290898
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 73368 273454 73688 273486
rect 73368 273218 73410 273454
rect 73646 273218 73688 273454
rect 73368 273134 73688 273218
rect 73368 272898 73410 273134
rect 73646 272898 73688 273134
rect 73368 272866 73688 272898
rect 104088 273454 104408 273486
rect 104088 273218 104130 273454
rect 104366 273218 104408 273454
rect 104088 273134 104408 273218
rect 104088 272898 104130 273134
rect 104366 272898 104408 273134
rect 104088 272866 104408 272898
rect 134808 273454 135128 273486
rect 134808 273218 134850 273454
rect 135086 273218 135128 273454
rect 134808 273134 135128 273218
rect 134808 272898 134850 273134
rect 135086 272898 135128 273134
rect 134808 272866 135128 272898
rect 165528 273454 165848 273486
rect 165528 273218 165570 273454
rect 165806 273218 165848 273454
rect 165528 273134 165848 273218
rect 165528 272898 165570 273134
rect 165806 272898 165848 273134
rect 165528 272866 165848 272898
rect 196248 273454 196568 273486
rect 196248 273218 196290 273454
rect 196526 273218 196568 273454
rect 196248 273134 196568 273218
rect 196248 272898 196290 273134
rect 196526 272898 196568 273134
rect 196248 272866 196568 272898
rect 226968 273454 227288 273486
rect 226968 273218 227010 273454
rect 227246 273218 227288 273454
rect 226968 273134 227288 273218
rect 226968 272898 227010 273134
rect 227246 272898 227288 273134
rect 226968 272866 227288 272898
rect 257688 273454 258008 273486
rect 257688 273218 257730 273454
rect 257966 273218 258008 273454
rect 257688 273134 258008 273218
rect 257688 272898 257730 273134
rect 257966 272898 258008 273134
rect 257688 272866 258008 272898
rect 288408 273454 288728 273486
rect 288408 273218 288450 273454
rect 288686 273218 288728 273454
rect 288408 273134 288728 273218
rect 288408 272898 288450 273134
rect 288686 272898 288728 273134
rect 288408 272866 288728 272898
rect 319128 273454 319448 273486
rect 319128 273218 319170 273454
rect 319406 273218 319448 273454
rect 319128 273134 319448 273218
rect 319128 272898 319170 273134
rect 319406 272898 319448 273134
rect 319128 272866 319448 272898
rect 349848 273454 350168 273486
rect 349848 273218 349890 273454
rect 350126 273218 350168 273454
rect 349848 273134 350168 273218
rect 349848 272898 349890 273134
rect 350126 272898 350168 273134
rect 349848 272866 350168 272898
rect 380568 273454 380888 273486
rect 380568 273218 380610 273454
rect 380846 273218 380888 273454
rect 380568 273134 380888 273218
rect 380568 272898 380610 273134
rect 380846 272898 380888 273134
rect 380568 272866 380888 272898
rect 411288 273454 411608 273486
rect 411288 273218 411330 273454
rect 411566 273218 411608 273454
rect 411288 273134 411608 273218
rect 411288 272898 411330 273134
rect 411566 272898 411608 273134
rect 411288 272866 411608 272898
rect 442008 273454 442328 273486
rect 442008 273218 442050 273454
rect 442286 273218 442328 273454
rect 442008 273134 442328 273218
rect 442008 272898 442050 273134
rect 442286 272898 442328 273134
rect 442008 272866 442328 272898
rect 472728 273454 473048 273486
rect 472728 273218 472770 273454
rect 473006 273218 473048 273454
rect 472728 273134 473048 273218
rect 472728 272898 472770 273134
rect 473006 272898 473048 273134
rect 472728 272866 473048 272898
rect 503448 273454 503768 273486
rect 503448 273218 503490 273454
rect 503726 273218 503768 273454
rect 503448 273134 503768 273218
rect 503448 272898 503490 273134
rect 503726 272898 503768 273134
rect 503448 272866 503768 272898
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 58008 255454 58328 255486
rect 58008 255218 58050 255454
rect 58286 255218 58328 255454
rect 58008 255134 58328 255218
rect 58008 254898 58050 255134
rect 58286 254898 58328 255134
rect 58008 254866 58328 254898
rect 88728 255454 89048 255486
rect 88728 255218 88770 255454
rect 89006 255218 89048 255454
rect 88728 255134 89048 255218
rect 88728 254898 88770 255134
rect 89006 254898 89048 255134
rect 88728 254866 89048 254898
rect 119448 255454 119768 255486
rect 119448 255218 119490 255454
rect 119726 255218 119768 255454
rect 119448 255134 119768 255218
rect 119448 254898 119490 255134
rect 119726 254898 119768 255134
rect 119448 254866 119768 254898
rect 150168 255454 150488 255486
rect 150168 255218 150210 255454
rect 150446 255218 150488 255454
rect 150168 255134 150488 255218
rect 150168 254898 150210 255134
rect 150446 254898 150488 255134
rect 150168 254866 150488 254898
rect 180888 255454 181208 255486
rect 180888 255218 180930 255454
rect 181166 255218 181208 255454
rect 180888 255134 181208 255218
rect 180888 254898 180930 255134
rect 181166 254898 181208 255134
rect 180888 254866 181208 254898
rect 211608 255454 211928 255486
rect 211608 255218 211650 255454
rect 211886 255218 211928 255454
rect 211608 255134 211928 255218
rect 211608 254898 211650 255134
rect 211886 254898 211928 255134
rect 211608 254866 211928 254898
rect 242328 255454 242648 255486
rect 242328 255218 242370 255454
rect 242606 255218 242648 255454
rect 242328 255134 242648 255218
rect 242328 254898 242370 255134
rect 242606 254898 242648 255134
rect 242328 254866 242648 254898
rect 273048 255454 273368 255486
rect 273048 255218 273090 255454
rect 273326 255218 273368 255454
rect 273048 255134 273368 255218
rect 273048 254898 273090 255134
rect 273326 254898 273368 255134
rect 273048 254866 273368 254898
rect 303768 255454 304088 255486
rect 303768 255218 303810 255454
rect 304046 255218 304088 255454
rect 303768 255134 304088 255218
rect 303768 254898 303810 255134
rect 304046 254898 304088 255134
rect 303768 254866 304088 254898
rect 334488 255454 334808 255486
rect 334488 255218 334530 255454
rect 334766 255218 334808 255454
rect 334488 255134 334808 255218
rect 334488 254898 334530 255134
rect 334766 254898 334808 255134
rect 334488 254866 334808 254898
rect 365208 255454 365528 255486
rect 365208 255218 365250 255454
rect 365486 255218 365528 255454
rect 365208 255134 365528 255218
rect 365208 254898 365250 255134
rect 365486 254898 365528 255134
rect 365208 254866 365528 254898
rect 395928 255454 396248 255486
rect 395928 255218 395970 255454
rect 396206 255218 396248 255454
rect 395928 255134 396248 255218
rect 395928 254898 395970 255134
rect 396206 254898 396248 255134
rect 395928 254866 396248 254898
rect 426648 255454 426968 255486
rect 426648 255218 426690 255454
rect 426926 255218 426968 255454
rect 426648 255134 426968 255218
rect 426648 254898 426690 255134
rect 426926 254898 426968 255134
rect 426648 254866 426968 254898
rect 457368 255454 457688 255486
rect 457368 255218 457410 255454
rect 457646 255218 457688 255454
rect 457368 255134 457688 255218
rect 457368 254898 457410 255134
rect 457646 254898 457688 255134
rect 457368 254866 457688 254898
rect 488088 255454 488408 255486
rect 488088 255218 488130 255454
rect 488366 255218 488408 255454
rect 488088 255134 488408 255218
rect 488088 254898 488130 255134
rect 488366 254898 488408 255134
rect 488088 254866 488408 254898
rect 518808 255454 519128 255486
rect 518808 255218 518850 255454
rect 519086 255218 519128 255454
rect 518808 255134 519128 255218
rect 518808 254898 518850 255134
rect 519086 254898 519128 255134
rect 518808 254866 519128 254898
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 73368 237454 73688 237486
rect 73368 237218 73410 237454
rect 73646 237218 73688 237454
rect 73368 237134 73688 237218
rect 73368 236898 73410 237134
rect 73646 236898 73688 237134
rect 73368 236866 73688 236898
rect 104088 237454 104408 237486
rect 104088 237218 104130 237454
rect 104366 237218 104408 237454
rect 104088 237134 104408 237218
rect 104088 236898 104130 237134
rect 104366 236898 104408 237134
rect 104088 236866 104408 236898
rect 134808 237454 135128 237486
rect 134808 237218 134850 237454
rect 135086 237218 135128 237454
rect 134808 237134 135128 237218
rect 134808 236898 134850 237134
rect 135086 236898 135128 237134
rect 134808 236866 135128 236898
rect 165528 237454 165848 237486
rect 165528 237218 165570 237454
rect 165806 237218 165848 237454
rect 165528 237134 165848 237218
rect 165528 236898 165570 237134
rect 165806 236898 165848 237134
rect 165528 236866 165848 236898
rect 196248 237454 196568 237486
rect 196248 237218 196290 237454
rect 196526 237218 196568 237454
rect 196248 237134 196568 237218
rect 196248 236898 196290 237134
rect 196526 236898 196568 237134
rect 196248 236866 196568 236898
rect 226968 237454 227288 237486
rect 226968 237218 227010 237454
rect 227246 237218 227288 237454
rect 226968 237134 227288 237218
rect 226968 236898 227010 237134
rect 227246 236898 227288 237134
rect 226968 236866 227288 236898
rect 257688 237454 258008 237486
rect 257688 237218 257730 237454
rect 257966 237218 258008 237454
rect 257688 237134 258008 237218
rect 257688 236898 257730 237134
rect 257966 236898 258008 237134
rect 257688 236866 258008 236898
rect 288408 237454 288728 237486
rect 288408 237218 288450 237454
rect 288686 237218 288728 237454
rect 288408 237134 288728 237218
rect 288408 236898 288450 237134
rect 288686 236898 288728 237134
rect 288408 236866 288728 236898
rect 319128 237454 319448 237486
rect 319128 237218 319170 237454
rect 319406 237218 319448 237454
rect 319128 237134 319448 237218
rect 319128 236898 319170 237134
rect 319406 236898 319448 237134
rect 319128 236866 319448 236898
rect 349848 237454 350168 237486
rect 349848 237218 349890 237454
rect 350126 237218 350168 237454
rect 349848 237134 350168 237218
rect 349848 236898 349890 237134
rect 350126 236898 350168 237134
rect 349848 236866 350168 236898
rect 380568 237454 380888 237486
rect 380568 237218 380610 237454
rect 380846 237218 380888 237454
rect 380568 237134 380888 237218
rect 380568 236898 380610 237134
rect 380846 236898 380888 237134
rect 380568 236866 380888 236898
rect 411288 237454 411608 237486
rect 411288 237218 411330 237454
rect 411566 237218 411608 237454
rect 411288 237134 411608 237218
rect 411288 236898 411330 237134
rect 411566 236898 411608 237134
rect 411288 236866 411608 236898
rect 442008 237454 442328 237486
rect 442008 237218 442050 237454
rect 442286 237218 442328 237454
rect 442008 237134 442328 237218
rect 442008 236898 442050 237134
rect 442286 236898 442328 237134
rect 442008 236866 442328 236898
rect 472728 237454 473048 237486
rect 472728 237218 472770 237454
rect 473006 237218 473048 237454
rect 472728 237134 473048 237218
rect 472728 236898 472770 237134
rect 473006 236898 473048 237134
rect 472728 236866 473048 236898
rect 503448 237454 503768 237486
rect 503448 237218 503490 237454
rect 503726 237218 503768 237454
rect 503448 237134 503768 237218
rect 503448 236898 503490 237134
rect 503726 236898 503768 237134
rect 503448 236866 503768 236898
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 58008 219454 58328 219486
rect 58008 219218 58050 219454
rect 58286 219218 58328 219454
rect 58008 219134 58328 219218
rect 58008 218898 58050 219134
rect 58286 218898 58328 219134
rect 58008 218866 58328 218898
rect 88728 219454 89048 219486
rect 88728 219218 88770 219454
rect 89006 219218 89048 219454
rect 88728 219134 89048 219218
rect 88728 218898 88770 219134
rect 89006 218898 89048 219134
rect 88728 218866 89048 218898
rect 119448 219454 119768 219486
rect 119448 219218 119490 219454
rect 119726 219218 119768 219454
rect 119448 219134 119768 219218
rect 119448 218898 119490 219134
rect 119726 218898 119768 219134
rect 119448 218866 119768 218898
rect 150168 219454 150488 219486
rect 150168 219218 150210 219454
rect 150446 219218 150488 219454
rect 150168 219134 150488 219218
rect 150168 218898 150210 219134
rect 150446 218898 150488 219134
rect 150168 218866 150488 218898
rect 180888 219454 181208 219486
rect 180888 219218 180930 219454
rect 181166 219218 181208 219454
rect 180888 219134 181208 219218
rect 180888 218898 180930 219134
rect 181166 218898 181208 219134
rect 180888 218866 181208 218898
rect 211608 219454 211928 219486
rect 211608 219218 211650 219454
rect 211886 219218 211928 219454
rect 211608 219134 211928 219218
rect 211608 218898 211650 219134
rect 211886 218898 211928 219134
rect 211608 218866 211928 218898
rect 242328 219454 242648 219486
rect 242328 219218 242370 219454
rect 242606 219218 242648 219454
rect 242328 219134 242648 219218
rect 242328 218898 242370 219134
rect 242606 218898 242648 219134
rect 242328 218866 242648 218898
rect 273048 219454 273368 219486
rect 273048 219218 273090 219454
rect 273326 219218 273368 219454
rect 273048 219134 273368 219218
rect 273048 218898 273090 219134
rect 273326 218898 273368 219134
rect 273048 218866 273368 218898
rect 303768 219454 304088 219486
rect 303768 219218 303810 219454
rect 304046 219218 304088 219454
rect 303768 219134 304088 219218
rect 303768 218898 303810 219134
rect 304046 218898 304088 219134
rect 303768 218866 304088 218898
rect 334488 219454 334808 219486
rect 334488 219218 334530 219454
rect 334766 219218 334808 219454
rect 334488 219134 334808 219218
rect 334488 218898 334530 219134
rect 334766 218898 334808 219134
rect 334488 218866 334808 218898
rect 365208 219454 365528 219486
rect 365208 219218 365250 219454
rect 365486 219218 365528 219454
rect 365208 219134 365528 219218
rect 365208 218898 365250 219134
rect 365486 218898 365528 219134
rect 365208 218866 365528 218898
rect 395928 219454 396248 219486
rect 395928 219218 395970 219454
rect 396206 219218 396248 219454
rect 395928 219134 396248 219218
rect 395928 218898 395970 219134
rect 396206 218898 396248 219134
rect 395928 218866 396248 218898
rect 426648 219454 426968 219486
rect 426648 219218 426690 219454
rect 426926 219218 426968 219454
rect 426648 219134 426968 219218
rect 426648 218898 426690 219134
rect 426926 218898 426968 219134
rect 426648 218866 426968 218898
rect 457368 219454 457688 219486
rect 457368 219218 457410 219454
rect 457646 219218 457688 219454
rect 457368 219134 457688 219218
rect 457368 218898 457410 219134
rect 457646 218898 457688 219134
rect 457368 218866 457688 218898
rect 488088 219454 488408 219486
rect 488088 219218 488130 219454
rect 488366 219218 488408 219454
rect 488088 219134 488408 219218
rect 488088 218898 488130 219134
rect 488366 218898 488408 219134
rect 488088 218866 488408 218898
rect 518808 219454 519128 219486
rect 518808 219218 518850 219454
rect 519086 219218 519128 219454
rect 518808 219134 519128 219218
rect 518808 218898 518850 219134
rect 519086 218898 519128 219134
rect 518808 218866 519128 218898
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 73368 201454 73688 201486
rect 73368 201218 73410 201454
rect 73646 201218 73688 201454
rect 73368 201134 73688 201218
rect 73368 200898 73410 201134
rect 73646 200898 73688 201134
rect 73368 200866 73688 200898
rect 104088 201454 104408 201486
rect 104088 201218 104130 201454
rect 104366 201218 104408 201454
rect 104088 201134 104408 201218
rect 104088 200898 104130 201134
rect 104366 200898 104408 201134
rect 104088 200866 104408 200898
rect 134808 201454 135128 201486
rect 134808 201218 134850 201454
rect 135086 201218 135128 201454
rect 134808 201134 135128 201218
rect 134808 200898 134850 201134
rect 135086 200898 135128 201134
rect 134808 200866 135128 200898
rect 165528 201454 165848 201486
rect 165528 201218 165570 201454
rect 165806 201218 165848 201454
rect 165528 201134 165848 201218
rect 165528 200898 165570 201134
rect 165806 200898 165848 201134
rect 165528 200866 165848 200898
rect 196248 201454 196568 201486
rect 196248 201218 196290 201454
rect 196526 201218 196568 201454
rect 196248 201134 196568 201218
rect 196248 200898 196290 201134
rect 196526 200898 196568 201134
rect 196248 200866 196568 200898
rect 226968 201454 227288 201486
rect 226968 201218 227010 201454
rect 227246 201218 227288 201454
rect 226968 201134 227288 201218
rect 226968 200898 227010 201134
rect 227246 200898 227288 201134
rect 226968 200866 227288 200898
rect 257688 201454 258008 201486
rect 257688 201218 257730 201454
rect 257966 201218 258008 201454
rect 257688 201134 258008 201218
rect 257688 200898 257730 201134
rect 257966 200898 258008 201134
rect 257688 200866 258008 200898
rect 288408 201454 288728 201486
rect 288408 201218 288450 201454
rect 288686 201218 288728 201454
rect 288408 201134 288728 201218
rect 288408 200898 288450 201134
rect 288686 200898 288728 201134
rect 288408 200866 288728 200898
rect 319128 201454 319448 201486
rect 319128 201218 319170 201454
rect 319406 201218 319448 201454
rect 319128 201134 319448 201218
rect 319128 200898 319170 201134
rect 319406 200898 319448 201134
rect 319128 200866 319448 200898
rect 349848 201454 350168 201486
rect 349848 201218 349890 201454
rect 350126 201218 350168 201454
rect 349848 201134 350168 201218
rect 349848 200898 349890 201134
rect 350126 200898 350168 201134
rect 349848 200866 350168 200898
rect 380568 201454 380888 201486
rect 380568 201218 380610 201454
rect 380846 201218 380888 201454
rect 380568 201134 380888 201218
rect 380568 200898 380610 201134
rect 380846 200898 380888 201134
rect 380568 200866 380888 200898
rect 411288 201454 411608 201486
rect 411288 201218 411330 201454
rect 411566 201218 411608 201454
rect 411288 201134 411608 201218
rect 411288 200898 411330 201134
rect 411566 200898 411608 201134
rect 411288 200866 411608 200898
rect 442008 201454 442328 201486
rect 442008 201218 442050 201454
rect 442286 201218 442328 201454
rect 442008 201134 442328 201218
rect 442008 200898 442050 201134
rect 442286 200898 442328 201134
rect 442008 200866 442328 200898
rect 472728 201454 473048 201486
rect 472728 201218 472770 201454
rect 473006 201218 473048 201454
rect 472728 201134 473048 201218
rect 472728 200898 472770 201134
rect 473006 200898 473048 201134
rect 472728 200866 473048 200898
rect 503448 201454 503768 201486
rect 503448 201218 503490 201454
rect 503726 201218 503768 201454
rect 503448 201134 503768 201218
rect 503448 200898 503490 201134
rect 503726 200898 503768 201134
rect 503448 200866 503768 200898
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 58008 183454 58328 183486
rect 58008 183218 58050 183454
rect 58286 183218 58328 183454
rect 58008 183134 58328 183218
rect 58008 182898 58050 183134
rect 58286 182898 58328 183134
rect 58008 182866 58328 182898
rect 88728 183454 89048 183486
rect 88728 183218 88770 183454
rect 89006 183218 89048 183454
rect 88728 183134 89048 183218
rect 88728 182898 88770 183134
rect 89006 182898 89048 183134
rect 88728 182866 89048 182898
rect 119448 183454 119768 183486
rect 119448 183218 119490 183454
rect 119726 183218 119768 183454
rect 119448 183134 119768 183218
rect 119448 182898 119490 183134
rect 119726 182898 119768 183134
rect 119448 182866 119768 182898
rect 150168 183454 150488 183486
rect 150168 183218 150210 183454
rect 150446 183218 150488 183454
rect 150168 183134 150488 183218
rect 150168 182898 150210 183134
rect 150446 182898 150488 183134
rect 150168 182866 150488 182898
rect 180888 183454 181208 183486
rect 180888 183218 180930 183454
rect 181166 183218 181208 183454
rect 180888 183134 181208 183218
rect 180888 182898 180930 183134
rect 181166 182898 181208 183134
rect 180888 182866 181208 182898
rect 211608 183454 211928 183486
rect 211608 183218 211650 183454
rect 211886 183218 211928 183454
rect 211608 183134 211928 183218
rect 211608 182898 211650 183134
rect 211886 182898 211928 183134
rect 211608 182866 211928 182898
rect 242328 183454 242648 183486
rect 242328 183218 242370 183454
rect 242606 183218 242648 183454
rect 242328 183134 242648 183218
rect 242328 182898 242370 183134
rect 242606 182898 242648 183134
rect 242328 182866 242648 182898
rect 273048 183454 273368 183486
rect 273048 183218 273090 183454
rect 273326 183218 273368 183454
rect 273048 183134 273368 183218
rect 273048 182898 273090 183134
rect 273326 182898 273368 183134
rect 273048 182866 273368 182898
rect 303768 183454 304088 183486
rect 303768 183218 303810 183454
rect 304046 183218 304088 183454
rect 303768 183134 304088 183218
rect 303768 182898 303810 183134
rect 304046 182898 304088 183134
rect 303768 182866 304088 182898
rect 334488 183454 334808 183486
rect 334488 183218 334530 183454
rect 334766 183218 334808 183454
rect 334488 183134 334808 183218
rect 334488 182898 334530 183134
rect 334766 182898 334808 183134
rect 334488 182866 334808 182898
rect 365208 183454 365528 183486
rect 365208 183218 365250 183454
rect 365486 183218 365528 183454
rect 365208 183134 365528 183218
rect 365208 182898 365250 183134
rect 365486 182898 365528 183134
rect 365208 182866 365528 182898
rect 395928 183454 396248 183486
rect 395928 183218 395970 183454
rect 396206 183218 396248 183454
rect 395928 183134 396248 183218
rect 395928 182898 395970 183134
rect 396206 182898 396248 183134
rect 395928 182866 396248 182898
rect 426648 183454 426968 183486
rect 426648 183218 426690 183454
rect 426926 183218 426968 183454
rect 426648 183134 426968 183218
rect 426648 182898 426690 183134
rect 426926 182898 426968 183134
rect 426648 182866 426968 182898
rect 457368 183454 457688 183486
rect 457368 183218 457410 183454
rect 457646 183218 457688 183454
rect 457368 183134 457688 183218
rect 457368 182898 457410 183134
rect 457646 182898 457688 183134
rect 457368 182866 457688 182898
rect 488088 183454 488408 183486
rect 488088 183218 488130 183454
rect 488366 183218 488408 183454
rect 488088 183134 488408 183218
rect 488088 182898 488130 183134
rect 488366 182898 488408 183134
rect 488088 182866 488408 182898
rect 518808 183454 519128 183486
rect 518808 183218 518850 183454
rect 519086 183218 519128 183454
rect 518808 183134 519128 183218
rect 518808 182898 518850 183134
rect 519086 182898 519128 183134
rect 518808 182866 519128 182898
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 73368 165454 73688 165486
rect 73368 165218 73410 165454
rect 73646 165218 73688 165454
rect 73368 165134 73688 165218
rect 73368 164898 73410 165134
rect 73646 164898 73688 165134
rect 73368 164866 73688 164898
rect 104088 165454 104408 165486
rect 104088 165218 104130 165454
rect 104366 165218 104408 165454
rect 104088 165134 104408 165218
rect 104088 164898 104130 165134
rect 104366 164898 104408 165134
rect 104088 164866 104408 164898
rect 134808 165454 135128 165486
rect 134808 165218 134850 165454
rect 135086 165218 135128 165454
rect 134808 165134 135128 165218
rect 134808 164898 134850 165134
rect 135086 164898 135128 165134
rect 134808 164866 135128 164898
rect 165528 165454 165848 165486
rect 165528 165218 165570 165454
rect 165806 165218 165848 165454
rect 165528 165134 165848 165218
rect 165528 164898 165570 165134
rect 165806 164898 165848 165134
rect 165528 164866 165848 164898
rect 196248 165454 196568 165486
rect 196248 165218 196290 165454
rect 196526 165218 196568 165454
rect 196248 165134 196568 165218
rect 196248 164898 196290 165134
rect 196526 164898 196568 165134
rect 196248 164866 196568 164898
rect 226968 165454 227288 165486
rect 226968 165218 227010 165454
rect 227246 165218 227288 165454
rect 226968 165134 227288 165218
rect 226968 164898 227010 165134
rect 227246 164898 227288 165134
rect 226968 164866 227288 164898
rect 257688 165454 258008 165486
rect 257688 165218 257730 165454
rect 257966 165218 258008 165454
rect 257688 165134 258008 165218
rect 257688 164898 257730 165134
rect 257966 164898 258008 165134
rect 257688 164866 258008 164898
rect 288408 165454 288728 165486
rect 288408 165218 288450 165454
rect 288686 165218 288728 165454
rect 288408 165134 288728 165218
rect 288408 164898 288450 165134
rect 288686 164898 288728 165134
rect 288408 164866 288728 164898
rect 319128 165454 319448 165486
rect 319128 165218 319170 165454
rect 319406 165218 319448 165454
rect 319128 165134 319448 165218
rect 319128 164898 319170 165134
rect 319406 164898 319448 165134
rect 319128 164866 319448 164898
rect 349848 165454 350168 165486
rect 349848 165218 349890 165454
rect 350126 165218 350168 165454
rect 349848 165134 350168 165218
rect 349848 164898 349890 165134
rect 350126 164898 350168 165134
rect 349848 164866 350168 164898
rect 380568 165454 380888 165486
rect 380568 165218 380610 165454
rect 380846 165218 380888 165454
rect 380568 165134 380888 165218
rect 380568 164898 380610 165134
rect 380846 164898 380888 165134
rect 380568 164866 380888 164898
rect 411288 165454 411608 165486
rect 411288 165218 411330 165454
rect 411566 165218 411608 165454
rect 411288 165134 411608 165218
rect 411288 164898 411330 165134
rect 411566 164898 411608 165134
rect 411288 164866 411608 164898
rect 442008 165454 442328 165486
rect 442008 165218 442050 165454
rect 442286 165218 442328 165454
rect 442008 165134 442328 165218
rect 442008 164898 442050 165134
rect 442286 164898 442328 165134
rect 442008 164866 442328 164898
rect 472728 165454 473048 165486
rect 472728 165218 472770 165454
rect 473006 165218 473048 165454
rect 472728 165134 473048 165218
rect 472728 164898 472770 165134
rect 473006 164898 473048 165134
rect 472728 164866 473048 164898
rect 503448 165454 503768 165486
rect 503448 165218 503490 165454
rect 503726 165218 503768 165454
rect 503448 165134 503768 165218
rect 503448 164898 503490 165134
rect 503726 164898 503768 165134
rect 503448 164866 503768 164898
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 58008 147454 58328 147486
rect 58008 147218 58050 147454
rect 58286 147218 58328 147454
rect 58008 147134 58328 147218
rect 58008 146898 58050 147134
rect 58286 146898 58328 147134
rect 58008 146866 58328 146898
rect 88728 147454 89048 147486
rect 88728 147218 88770 147454
rect 89006 147218 89048 147454
rect 88728 147134 89048 147218
rect 88728 146898 88770 147134
rect 89006 146898 89048 147134
rect 88728 146866 89048 146898
rect 119448 147454 119768 147486
rect 119448 147218 119490 147454
rect 119726 147218 119768 147454
rect 119448 147134 119768 147218
rect 119448 146898 119490 147134
rect 119726 146898 119768 147134
rect 119448 146866 119768 146898
rect 150168 147454 150488 147486
rect 150168 147218 150210 147454
rect 150446 147218 150488 147454
rect 150168 147134 150488 147218
rect 150168 146898 150210 147134
rect 150446 146898 150488 147134
rect 150168 146866 150488 146898
rect 180888 147454 181208 147486
rect 180888 147218 180930 147454
rect 181166 147218 181208 147454
rect 180888 147134 181208 147218
rect 180888 146898 180930 147134
rect 181166 146898 181208 147134
rect 180888 146866 181208 146898
rect 211608 147454 211928 147486
rect 211608 147218 211650 147454
rect 211886 147218 211928 147454
rect 211608 147134 211928 147218
rect 211608 146898 211650 147134
rect 211886 146898 211928 147134
rect 211608 146866 211928 146898
rect 242328 147454 242648 147486
rect 242328 147218 242370 147454
rect 242606 147218 242648 147454
rect 242328 147134 242648 147218
rect 242328 146898 242370 147134
rect 242606 146898 242648 147134
rect 242328 146866 242648 146898
rect 273048 147454 273368 147486
rect 273048 147218 273090 147454
rect 273326 147218 273368 147454
rect 273048 147134 273368 147218
rect 273048 146898 273090 147134
rect 273326 146898 273368 147134
rect 273048 146866 273368 146898
rect 303768 147454 304088 147486
rect 303768 147218 303810 147454
rect 304046 147218 304088 147454
rect 303768 147134 304088 147218
rect 303768 146898 303810 147134
rect 304046 146898 304088 147134
rect 303768 146866 304088 146898
rect 334488 147454 334808 147486
rect 334488 147218 334530 147454
rect 334766 147218 334808 147454
rect 334488 147134 334808 147218
rect 334488 146898 334530 147134
rect 334766 146898 334808 147134
rect 334488 146866 334808 146898
rect 365208 147454 365528 147486
rect 365208 147218 365250 147454
rect 365486 147218 365528 147454
rect 365208 147134 365528 147218
rect 365208 146898 365250 147134
rect 365486 146898 365528 147134
rect 365208 146866 365528 146898
rect 395928 147454 396248 147486
rect 395928 147218 395970 147454
rect 396206 147218 396248 147454
rect 395928 147134 396248 147218
rect 395928 146898 395970 147134
rect 396206 146898 396248 147134
rect 395928 146866 396248 146898
rect 426648 147454 426968 147486
rect 426648 147218 426690 147454
rect 426926 147218 426968 147454
rect 426648 147134 426968 147218
rect 426648 146898 426690 147134
rect 426926 146898 426968 147134
rect 426648 146866 426968 146898
rect 457368 147454 457688 147486
rect 457368 147218 457410 147454
rect 457646 147218 457688 147454
rect 457368 147134 457688 147218
rect 457368 146898 457410 147134
rect 457646 146898 457688 147134
rect 457368 146866 457688 146898
rect 488088 147454 488408 147486
rect 488088 147218 488130 147454
rect 488366 147218 488408 147454
rect 488088 147134 488408 147218
rect 488088 146898 488130 147134
rect 488366 146898 488408 147134
rect 488088 146866 488408 146898
rect 518808 147454 519128 147486
rect 518808 147218 518850 147454
rect 519086 147218 519128 147454
rect 518808 147134 519128 147218
rect 518808 146898 518850 147134
rect 519086 146898 519128 147134
rect 518808 146866 519128 146898
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 73368 129454 73688 129486
rect 73368 129218 73410 129454
rect 73646 129218 73688 129454
rect 73368 129134 73688 129218
rect 73368 128898 73410 129134
rect 73646 128898 73688 129134
rect 73368 128866 73688 128898
rect 104088 129454 104408 129486
rect 104088 129218 104130 129454
rect 104366 129218 104408 129454
rect 104088 129134 104408 129218
rect 104088 128898 104130 129134
rect 104366 128898 104408 129134
rect 104088 128866 104408 128898
rect 134808 129454 135128 129486
rect 134808 129218 134850 129454
rect 135086 129218 135128 129454
rect 134808 129134 135128 129218
rect 134808 128898 134850 129134
rect 135086 128898 135128 129134
rect 134808 128866 135128 128898
rect 165528 129454 165848 129486
rect 165528 129218 165570 129454
rect 165806 129218 165848 129454
rect 165528 129134 165848 129218
rect 165528 128898 165570 129134
rect 165806 128898 165848 129134
rect 165528 128866 165848 128898
rect 196248 129454 196568 129486
rect 196248 129218 196290 129454
rect 196526 129218 196568 129454
rect 196248 129134 196568 129218
rect 196248 128898 196290 129134
rect 196526 128898 196568 129134
rect 196248 128866 196568 128898
rect 226968 129454 227288 129486
rect 226968 129218 227010 129454
rect 227246 129218 227288 129454
rect 226968 129134 227288 129218
rect 226968 128898 227010 129134
rect 227246 128898 227288 129134
rect 226968 128866 227288 128898
rect 257688 129454 258008 129486
rect 257688 129218 257730 129454
rect 257966 129218 258008 129454
rect 257688 129134 258008 129218
rect 257688 128898 257730 129134
rect 257966 128898 258008 129134
rect 257688 128866 258008 128898
rect 288408 129454 288728 129486
rect 288408 129218 288450 129454
rect 288686 129218 288728 129454
rect 288408 129134 288728 129218
rect 288408 128898 288450 129134
rect 288686 128898 288728 129134
rect 288408 128866 288728 128898
rect 319128 129454 319448 129486
rect 319128 129218 319170 129454
rect 319406 129218 319448 129454
rect 319128 129134 319448 129218
rect 319128 128898 319170 129134
rect 319406 128898 319448 129134
rect 319128 128866 319448 128898
rect 349848 129454 350168 129486
rect 349848 129218 349890 129454
rect 350126 129218 350168 129454
rect 349848 129134 350168 129218
rect 349848 128898 349890 129134
rect 350126 128898 350168 129134
rect 349848 128866 350168 128898
rect 380568 129454 380888 129486
rect 380568 129218 380610 129454
rect 380846 129218 380888 129454
rect 380568 129134 380888 129218
rect 380568 128898 380610 129134
rect 380846 128898 380888 129134
rect 380568 128866 380888 128898
rect 411288 129454 411608 129486
rect 411288 129218 411330 129454
rect 411566 129218 411608 129454
rect 411288 129134 411608 129218
rect 411288 128898 411330 129134
rect 411566 128898 411608 129134
rect 411288 128866 411608 128898
rect 442008 129454 442328 129486
rect 442008 129218 442050 129454
rect 442286 129218 442328 129454
rect 442008 129134 442328 129218
rect 442008 128898 442050 129134
rect 442286 128898 442328 129134
rect 442008 128866 442328 128898
rect 472728 129454 473048 129486
rect 472728 129218 472770 129454
rect 473006 129218 473048 129454
rect 472728 129134 473048 129218
rect 472728 128898 472770 129134
rect 473006 128898 473048 129134
rect 472728 128866 473048 128898
rect 503448 129454 503768 129486
rect 503448 129218 503490 129454
rect 503726 129218 503768 129454
rect 503448 129134 503768 129218
rect 503448 128898 503490 129134
rect 503726 128898 503768 129134
rect 503448 128866 503768 128898
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 58008 111454 58328 111486
rect 58008 111218 58050 111454
rect 58286 111218 58328 111454
rect 58008 111134 58328 111218
rect 58008 110898 58050 111134
rect 58286 110898 58328 111134
rect 58008 110866 58328 110898
rect 88728 111454 89048 111486
rect 88728 111218 88770 111454
rect 89006 111218 89048 111454
rect 88728 111134 89048 111218
rect 88728 110898 88770 111134
rect 89006 110898 89048 111134
rect 88728 110866 89048 110898
rect 119448 111454 119768 111486
rect 119448 111218 119490 111454
rect 119726 111218 119768 111454
rect 119448 111134 119768 111218
rect 119448 110898 119490 111134
rect 119726 110898 119768 111134
rect 119448 110866 119768 110898
rect 150168 111454 150488 111486
rect 150168 111218 150210 111454
rect 150446 111218 150488 111454
rect 150168 111134 150488 111218
rect 150168 110898 150210 111134
rect 150446 110898 150488 111134
rect 150168 110866 150488 110898
rect 180888 111454 181208 111486
rect 180888 111218 180930 111454
rect 181166 111218 181208 111454
rect 180888 111134 181208 111218
rect 180888 110898 180930 111134
rect 181166 110898 181208 111134
rect 180888 110866 181208 110898
rect 211608 111454 211928 111486
rect 211608 111218 211650 111454
rect 211886 111218 211928 111454
rect 211608 111134 211928 111218
rect 211608 110898 211650 111134
rect 211886 110898 211928 111134
rect 211608 110866 211928 110898
rect 242328 111454 242648 111486
rect 242328 111218 242370 111454
rect 242606 111218 242648 111454
rect 242328 111134 242648 111218
rect 242328 110898 242370 111134
rect 242606 110898 242648 111134
rect 242328 110866 242648 110898
rect 273048 111454 273368 111486
rect 273048 111218 273090 111454
rect 273326 111218 273368 111454
rect 273048 111134 273368 111218
rect 273048 110898 273090 111134
rect 273326 110898 273368 111134
rect 273048 110866 273368 110898
rect 303768 111454 304088 111486
rect 303768 111218 303810 111454
rect 304046 111218 304088 111454
rect 303768 111134 304088 111218
rect 303768 110898 303810 111134
rect 304046 110898 304088 111134
rect 303768 110866 304088 110898
rect 334488 111454 334808 111486
rect 334488 111218 334530 111454
rect 334766 111218 334808 111454
rect 334488 111134 334808 111218
rect 334488 110898 334530 111134
rect 334766 110898 334808 111134
rect 334488 110866 334808 110898
rect 365208 111454 365528 111486
rect 365208 111218 365250 111454
rect 365486 111218 365528 111454
rect 365208 111134 365528 111218
rect 365208 110898 365250 111134
rect 365486 110898 365528 111134
rect 365208 110866 365528 110898
rect 395928 111454 396248 111486
rect 395928 111218 395970 111454
rect 396206 111218 396248 111454
rect 395928 111134 396248 111218
rect 395928 110898 395970 111134
rect 396206 110898 396248 111134
rect 395928 110866 396248 110898
rect 426648 111454 426968 111486
rect 426648 111218 426690 111454
rect 426926 111218 426968 111454
rect 426648 111134 426968 111218
rect 426648 110898 426690 111134
rect 426926 110898 426968 111134
rect 426648 110866 426968 110898
rect 457368 111454 457688 111486
rect 457368 111218 457410 111454
rect 457646 111218 457688 111454
rect 457368 111134 457688 111218
rect 457368 110898 457410 111134
rect 457646 110898 457688 111134
rect 457368 110866 457688 110898
rect 488088 111454 488408 111486
rect 488088 111218 488130 111454
rect 488366 111218 488408 111454
rect 488088 111134 488408 111218
rect 488088 110898 488130 111134
rect 488366 110898 488408 111134
rect 488088 110866 488408 110898
rect 518808 111454 519128 111486
rect 518808 111218 518850 111454
rect 519086 111218 519128 111454
rect 518808 111134 519128 111218
rect 518808 110898 518850 111134
rect 519086 110898 519128 111134
rect 518808 110866 519128 110898
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 73368 93454 73688 93486
rect 73368 93218 73410 93454
rect 73646 93218 73688 93454
rect 73368 93134 73688 93218
rect 73368 92898 73410 93134
rect 73646 92898 73688 93134
rect 73368 92866 73688 92898
rect 104088 93454 104408 93486
rect 104088 93218 104130 93454
rect 104366 93218 104408 93454
rect 104088 93134 104408 93218
rect 104088 92898 104130 93134
rect 104366 92898 104408 93134
rect 104088 92866 104408 92898
rect 134808 93454 135128 93486
rect 134808 93218 134850 93454
rect 135086 93218 135128 93454
rect 134808 93134 135128 93218
rect 134808 92898 134850 93134
rect 135086 92898 135128 93134
rect 134808 92866 135128 92898
rect 165528 93454 165848 93486
rect 165528 93218 165570 93454
rect 165806 93218 165848 93454
rect 165528 93134 165848 93218
rect 165528 92898 165570 93134
rect 165806 92898 165848 93134
rect 165528 92866 165848 92898
rect 196248 93454 196568 93486
rect 196248 93218 196290 93454
rect 196526 93218 196568 93454
rect 196248 93134 196568 93218
rect 196248 92898 196290 93134
rect 196526 92898 196568 93134
rect 196248 92866 196568 92898
rect 226968 93454 227288 93486
rect 226968 93218 227010 93454
rect 227246 93218 227288 93454
rect 226968 93134 227288 93218
rect 226968 92898 227010 93134
rect 227246 92898 227288 93134
rect 226968 92866 227288 92898
rect 257688 93454 258008 93486
rect 257688 93218 257730 93454
rect 257966 93218 258008 93454
rect 257688 93134 258008 93218
rect 257688 92898 257730 93134
rect 257966 92898 258008 93134
rect 257688 92866 258008 92898
rect 288408 93454 288728 93486
rect 288408 93218 288450 93454
rect 288686 93218 288728 93454
rect 288408 93134 288728 93218
rect 288408 92898 288450 93134
rect 288686 92898 288728 93134
rect 288408 92866 288728 92898
rect 319128 93454 319448 93486
rect 319128 93218 319170 93454
rect 319406 93218 319448 93454
rect 319128 93134 319448 93218
rect 319128 92898 319170 93134
rect 319406 92898 319448 93134
rect 319128 92866 319448 92898
rect 349848 93454 350168 93486
rect 349848 93218 349890 93454
rect 350126 93218 350168 93454
rect 349848 93134 350168 93218
rect 349848 92898 349890 93134
rect 350126 92898 350168 93134
rect 349848 92866 350168 92898
rect 380568 93454 380888 93486
rect 380568 93218 380610 93454
rect 380846 93218 380888 93454
rect 380568 93134 380888 93218
rect 380568 92898 380610 93134
rect 380846 92898 380888 93134
rect 380568 92866 380888 92898
rect 411288 93454 411608 93486
rect 411288 93218 411330 93454
rect 411566 93218 411608 93454
rect 411288 93134 411608 93218
rect 411288 92898 411330 93134
rect 411566 92898 411608 93134
rect 411288 92866 411608 92898
rect 442008 93454 442328 93486
rect 442008 93218 442050 93454
rect 442286 93218 442328 93454
rect 442008 93134 442328 93218
rect 442008 92898 442050 93134
rect 442286 92898 442328 93134
rect 442008 92866 442328 92898
rect 472728 93454 473048 93486
rect 472728 93218 472770 93454
rect 473006 93218 473048 93454
rect 472728 93134 473048 93218
rect 472728 92898 472770 93134
rect 473006 92898 473048 93134
rect 472728 92866 473048 92898
rect 503448 93454 503768 93486
rect 503448 93218 503490 93454
rect 503726 93218 503768 93454
rect 503448 93134 503768 93218
rect 503448 92898 503490 93134
rect 503726 92898 503768 93134
rect 503448 92866 503768 92898
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 58008 75454 58328 75486
rect 58008 75218 58050 75454
rect 58286 75218 58328 75454
rect 58008 75134 58328 75218
rect 58008 74898 58050 75134
rect 58286 74898 58328 75134
rect 58008 74866 58328 74898
rect 88728 75454 89048 75486
rect 88728 75218 88770 75454
rect 89006 75218 89048 75454
rect 88728 75134 89048 75218
rect 88728 74898 88770 75134
rect 89006 74898 89048 75134
rect 88728 74866 89048 74898
rect 119448 75454 119768 75486
rect 119448 75218 119490 75454
rect 119726 75218 119768 75454
rect 119448 75134 119768 75218
rect 119448 74898 119490 75134
rect 119726 74898 119768 75134
rect 119448 74866 119768 74898
rect 150168 75454 150488 75486
rect 150168 75218 150210 75454
rect 150446 75218 150488 75454
rect 150168 75134 150488 75218
rect 150168 74898 150210 75134
rect 150446 74898 150488 75134
rect 150168 74866 150488 74898
rect 180888 75454 181208 75486
rect 180888 75218 180930 75454
rect 181166 75218 181208 75454
rect 180888 75134 181208 75218
rect 180888 74898 180930 75134
rect 181166 74898 181208 75134
rect 180888 74866 181208 74898
rect 211608 75454 211928 75486
rect 211608 75218 211650 75454
rect 211886 75218 211928 75454
rect 211608 75134 211928 75218
rect 211608 74898 211650 75134
rect 211886 74898 211928 75134
rect 211608 74866 211928 74898
rect 242328 75454 242648 75486
rect 242328 75218 242370 75454
rect 242606 75218 242648 75454
rect 242328 75134 242648 75218
rect 242328 74898 242370 75134
rect 242606 74898 242648 75134
rect 242328 74866 242648 74898
rect 273048 75454 273368 75486
rect 273048 75218 273090 75454
rect 273326 75218 273368 75454
rect 273048 75134 273368 75218
rect 273048 74898 273090 75134
rect 273326 74898 273368 75134
rect 273048 74866 273368 74898
rect 303768 75454 304088 75486
rect 303768 75218 303810 75454
rect 304046 75218 304088 75454
rect 303768 75134 304088 75218
rect 303768 74898 303810 75134
rect 304046 74898 304088 75134
rect 303768 74866 304088 74898
rect 334488 75454 334808 75486
rect 334488 75218 334530 75454
rect 334766 75218 334808 75454
rect 334488 75134 334808 75218
rect 334488 74898 334530 75134
rect 334766 74898 334808 75134
rect 334488 74866 334808 74898
rect 365208 75454 365528 75486
rect 365208 75218 365250 75454
rect 365486 75218 365528 75454
rect 365208 75134 365528 75218
rect 365208 74898 365250 75134
rect 365486 74898 365528 75134
rect 365208 74866 365528 74898
rect 395928 75454 396248 75486
rect 395928 75218 395970 75454
rect 396206 75218 396248 75454
rect 395928 75134 396248 75218
rect 395928 74898 395970 75134
rect 396206 74898 396248 75134
rect 395928 74866 396248 74898
rect 426648 75454 426968 75486
rect 426648 75218 426690 75454
rect 426926 75218 426968 75454
rect 426648 75134 426968 75218
rect 426648 74898 426690 75134
rect 426926 74898 426968 75134
rect 426648 74866 426968 74898
rect 457368 75454 457688 75486
rect 457368 75218 457410 75454
rect 457646 75218 457688 75454
rect 457368 75134 457688 75218
rect 457368 74898 457410 75134
rect 457646 74898 457688 75134
rect 457368 74866 457688 74898
rect 488088 75454 488408 75486
rect 488088 75218 488130 75454
rect 488366 75218 488408 75454
rect 488088 75134 488408 75218
rect 488088 74898 488130 75134
rect 488366 74898 488408 75134
rect 488088 74866 488408 74898
rect 518808 75454 519128 75486
rect 518808 75218 518850 75454
rect 519086 75218 519128 75454
rect 518808 75134 519128 75218
rect 518808 74898 518850 75134
rect 519086 74898 519128 75134
rect 518808 74866 519128 74898
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 57454 56414 63400
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 61174 60134 63400
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 63400
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 63400
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 63400
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 63400
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 63400
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 63400
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 63400
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 63400
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 63400
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 63400
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 63400
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 63400
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 63400
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 63400
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 63400
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 63400
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 63400
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 63400
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 63400
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 63400
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 63400
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 63400
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 63400
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 63400
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 63400
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 63400
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 63400
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 63400
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 63400
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 63400
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 63400
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 63400
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 63400
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 63400
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 63400
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 63400
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 63400
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 63400
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 63400
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 63400
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 63400
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 63400
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 63400
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 63400
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 63400
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 63400
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 63400
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 63400
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 63400
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 63400
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 63400
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 63400
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 63400
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 63400
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 63400
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 63400
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 63400
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 63400
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 63400
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 63400
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 63400
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 63400
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 63400
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 61174 348134 63400
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 63400
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 63400
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 63400
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 63400
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 63400
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 63400
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 63400
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 61174 384134 63400
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 63400
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 63400
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 63400
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 63400
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 63400
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 63400
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 63400
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 61174 420134 63400
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 63400
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 63400
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 63400
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 63400
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 63400
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 63400
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 63400
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 61174 456134 63400
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 63400
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 63400
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 63400
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 63400
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 63400
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 63400
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 63400
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 61174 492134 63400
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 63400
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 63400
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 63400
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 63400
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 63400
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 63400
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 63400
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 61174 528134 63400
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 63400
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 73410 633218 73646 633454
rect 73410 632898 73646 633134
rect 104130 633218 104366 633454
rect 104130 632898 104366 633134
rect 134850 633218 135086 633454
rect 134850 632898 135086 633134
rect 165570 633218 165806 633454
rect 165570 632898 165806 633134
rect 196290 633218 196526 633454
rect 196290 632898 196526 633134
rect 227010 633218 227246 633454
rect 227010 632898 227246 633134
rect 257730 633218 257966 633454
rect 257730 632898 257966 633134
rect 288450 633218 288686 633454
rect 288450 632898 288686 633134
rect 319170 633218 319406 633454
rect 319170 632898 319406 633134
rect 349890 633218 350126 633454
rect 349890 632898 350126 633134
rect 380610 633218 380846 633454
rect 380610 632898 380846 633134
rect 411330 633218 411566 633454
rect 411330 632898 411566 633134
rect 442050 633218 442286 633454
rect 442050 632898 442286 633134
rect 472770 633218 473006 633454
rect 472770 632898 473006 633134
rect 503490 633218 503726 633454
rect 503490 632898 503726 633134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 58050 615218 58286 615454
rect 58050 614898 58286 615134
rect 88770 615218 89006 615454
rect 88770 614898 89006 615134
rect 119490 615218 119726 615454
rect 119490 614898 119726 615134
rect 150210 615218 150446 615454
rect 150210 614898 150446 615134
rect 180930 615218 181166 615454
rect 180930 614898 181166 615134
rect 211650 615218 211886 615454
rect 211650 614898 211886 615134
rect 242370 615218 242606 615454
rect 242370 614898 242606 615134
rect 273090 615218 273326 615454
rect 273090 614898 273326 615134
rect 303810 615218 304046 615454
rect 303810 614898 304046 615134
rect 334530 615218 334766 615454
rect 334530 614898 334766 615134
rect 365250 615218 365486 615454
rect 365250 614898 365486 615134
rect 395970 615218 396206 615454
rect 395970 614898 396206 615134
rect 426690 615218 426926 615454
rect 426690 614898 426926 615134
rect 457410 615218 457646 615454
rect 457410 614898 457646 615134
rect 488130 615218 488366 615454
rect 488130 614898 488366 615134
rect 518850 615218 519086 615454
rect 518850 614898 519086 615134
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 73410 597218 73646 597454
rect 73410 596898 73646 597134
rect 104130 597218 104366 597454
rect 104130 596898 104366 597134
rect 134850 597218 135086 597454
rect 134850 596898 135086 597134
rect 165570 597218 165806 597454
rect 165570 596898 165806 597134
rect 196290 597218 196526 597454
rect 196290 596898 196526 597134
rect 227010 597218 227246 597454
rect 227010 596898 227246 597134
rect 257730 597218 257966 597454
rect 257730 596898 257966 597134
rect 288450 597218 288686 597454
rect 288450 596898 288686 597134
rect 319170 597218 319406 597454
rect 319170 596898 319406 597134
rect 349890 597218 350126 597454
rect 349890 596898 350126 597134
rect 380610 597218 380846 597454
rect 380610 596898 380846 597134
rect 411330 597218 411566 597454
rect 411330 596898 411566 597134
rect 442050 597218 442286 597454
rect 442050 596898 442286 597134
rect 472770 597218 473006 597454
rect 472770 596898 473006 597134
rect 503490 597218 503726 597454
rect 503490 596898 503726 597134
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 58050 579218 58286 579454
rect 58050 578898 58286 579134
rect 88770 579218 89006 579454
rect 88770 578898 89006 579134
rect 119490 579218 119726 579454
rect 119490 578898 119726 579134
rect 150210 579218 150446 579454
rect 150210 578898 150446 579134
rect 180930 579218 181166 579454
rect 180930 578898 181166 579134
rect 211650 579218 211886 579454
rect 211650 578898 211886 579134
rect 242370 579218 242606 579454
rect 242370 578898 242606 579134
rect 273090 579218 273326 579454
rect 273090 578898 273326 579134
rect 303810 579218 304046 579454
rect 303810 578898 304046 579134
rect 334530 579218 334766 579454
rect 334530 578898 334766 579134
rect 365250 579218 365486 579454
rect 365250 578898 365486 579134
rect 395970 579218 396206 579454
rect 395970 578898 396206 579134
rect 426690 579218 426926 579454
rect 426690 578898 426926 579134
rect 457410 579218 457646 579454
rect 457410 578898 457646 579134
rect 488130 579218 488366 579454
rect 488130 578898 488366 579134
rect 518850 579218 519086 579454
rect 518850 578898 519086 579134
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 73410 561218 73646 561454
rect 73410 560898 73646 561134
rect 104130 561218 104366 561454
rect 104130 560898 104366 561134
rect 134850 561218 135086 561454
rect 134850 560898 135086 561134
rect 165570 561218 165806 561454
rect 165570 560898 165806 561134
rect 196290 561218 196526 561454
rect 196290 560898 196526 561134
rect 227010 561218 227246 561454
rect 227010 560898 227246 561134
rect 257730 561218 257966 561454
rect 257730 560898 257966 561134
rect 288450 561218 288686 561454
rect 288450 560898 288686 561134
rect 319170 561218 319406 561454
rect 319170 560898 319406 561134
rect 349890 561218 350126 561454
rect 349890 560898 350126 561134
rect 380610 561218 380846 561454
rect 380610 560898 380846 561134
rect 411330 561218 411566 561454
rect 411330 560898 411566 561134
rect 442050 561218 442286 561454
rect 442050 560898 442286 561134
rect 472770 561218 473006 561454
rect 472770 560898 473006 561134
rect 503490 561218 503726 561454
rect 503490 560898 503726 561134
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 58050 543218 58286 543454
rect 58050 542898 58286 543134
rect 88770 543218 89006 543454
rect 88770 542898 89006 543134
rect 119490 543218 119726 543454
rect 119490 542898 119726 543134
rect 150210 543218 150446 543454
rect 150210 542898 150446 543134
rect 180930 543218 181166 543454
rect 180930 542898 181166 543134
rect 211650 543218 211886 543454
rect 211650 542898 211886 543134
rect 242370 543218 242606 543454
rect 242370 542898 242606 543134
rect 273090 543218 273326 543454
rect 273090 542898 273326 543134
rect 303810 543218 304046 543454
rect 303810 542898 304046 543134
rect 334530 543218 334766 543454
rect 334530 542898 334766 543134
rect 365250 543218 365486 543454
rect 365250 542898 365486 543134
rect 395970 543218 396206 543454
rect 395970 542898 396206 543134
rect 426690 543218 426926 543454
rect 426690 542898 426926 543134
rect 457410 543218 457646 543454
rect 457410 542898 457646 543134
rect 488130 543218 488366 543454
rect 488130 542898 488366 543134
rect 518850 543218 519086 543454
rect 518850 542898 519086 543134
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 73410 525218 73646 525454
rect 73410 524898 73646 525134
rect 104130 525218 104366 525454
rect 104130 524898 104366 525134
rect 134850 525218 135086 525454
rect 134850 524898 135086 525134
rect 165570 525218 165806 525454
rect 165570 524898 165806 525134
rect 196290 525218 196526 525454
rect 196290 524898 196526 525134
rect 227010 525218 227246 525454
rect 227010 524898 227246 525134
rect 257730 525218 257966 525454
rect 257730 524898 257966 525134
rect 288450 525218 288686 525454
rect 288450 524898 288686 525134
rect 319170 525218 319406 525454
rect 319170 524898 319406 525134
rect 349890 525218 350126 525454
rect 349890 524898 350126 525134
rect 380610 525218 380846 525454
rect 380610 524898 380846 525134
rect 411330 525218 411566 525454
rect 411330 524898 411566 525134
rect 442050 525218 442286 525454
rect 442050 524898 442286 525134
rect 472770 525218 473006 525454
rect 472770 524898 473006 525134
rect 503490 525218 503726 525454
rect 503490 524898 503726 525134
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 58050 507218 58286 507454
rect 58050 506898 58286 507134
rect 88770 507218 89006 507454
rect 88770 506898 89006 507134
rect 119490 507218 119726 507454
rect 119490 506898 119726 507134
rect 150210 507218 150446 507454
rect 150210 506898 150446 507134
rect 180930 507218 181166 507454
rect 180930 506898 181166 507134
rect 211650 507218 211886 507454
rect 211650 506898 211886 507134
rect 242370 507218 242606 507454
rect 242370 506898 242606 507134
rect 273090 507218 273326 507454
rect 273090 506898 273326 507134
rect 303810 507218 304046 507454
rect 303810 506898 304046 507134
rect 334530 507218 334766 507454
rect 334530 506898 334766 507134
rect 365250 507218 365486 507454
rect 365250 506898 365486 507134
rect 395970 507218 396206 507454
rect 395970 506898 396206 507134
rect 426690 507218 426926 507454
rect 426690 506898 426926 507134
rect 457410 507218 457646 507454
rect 457410 506898 457646 507134
rect 488130 507218 488366 507454
rect 488130 506898 488366 507134
rect 518850 507218 519086 507454
rect 518850 506898 519086 507134
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 73410 489218 73646 489454
rect 73410 488898 73646 489134
rect 104130 489218 104366 489454
rect 104130 488898 104366 489134
rect 134850 489218 135086 489454
rect 134850 488898 135086 489134
rect 165570 489218 165806 489454
rect 165570 488898 165806 489134
rect 196290 489218 196526 489454
rect 196290 488898 196526 489134
rect 227010 489218 227246 489454
rect 227010 488898 227246 489134
rect 257730 489218 257966 489454
rect 257730 488898 257966 489134
rect 288450 489218 288686 489454
rect 288450 488898 288686 489134
rect 319170 489218 319406 489454
rect 319170 488898 319406 489134
rect 349890 489218 350126 489454
rect 349890 488898 350126 489134
rect 380610 489218 380846 489454
rect 380610 488898 380846 489134
rect 411330 489218 411566 489454
rect 411330 488898 411566 489134
rect 442050 489218 442286 489454
rect 442050 488898 442286 489134
rect 472770 489218 473006 489454
rect 472770 488898 473006 489134
rect 503490 489218 503726 489454
rect 503490 488898 503726 489134
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 58050 471218 58286 471454
rect 58050 470898 58286 471134
rect 88770 471218 89006 471454
rect 88770 470898 89006 471134
rect 119490 471218 119726 471454
rect 119490 470898 119726 471134
rect 150210 471218 150446 471454
rect 150210 470898 150446 471134
rect 180930 471218 181166 471454
rect 180930 470898 181166 471134
rect 211650 471218 211886 471454
rect 211650 470898 211886 471134
rect 242370 471218 242606 471454
rect 242370 470898 242606 471134
rect 273090 471218 273326 471454
rect 273090 470898 273326 471134
rect 303810 471218 304046 471454
rect 303810 470898 304046 471134
rect 334530 471218 334766 471454
rect 334530 470898 334766 471134
rect 365250 471218 365486 471454
rect 365250 470898 365486 471134
rect 395970 471218 396206 471454
rect 395970 470898 396206 471134
rect 426690 471218 426926 471454
rect 426690 470898 426926 471134
rect 457410 471218 457646 471454
rect 457410 470898 457646 471134
rect 488130 471218 488366 471454
rect 488130 470898 488366 471134
rect 518850 471218 519086 471454
rect 518850 470898 519086 471134
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 73410 453218 73646 453454
rect 73410 452898 73646 453134
rect 104130 453218 104366 453454
rect 104130 452898 104366 453134
rect 134850 453218 135086 453454
rect 134850 452898 135086 453134
rect 165570 453218 165806 453454
rect 165570 452898 165806 453134
rect 196290 453218 196526 453454
rect 196290 452898 196526 453134
rect 227010 453218 227246 453454
rect 227010 452898 227246 453134
rect 257730 453218 257966 453454
rect 257730 452898 257966 453134
rect 288450 453218 288686 453454
rect 288450 452898 288686 453134
rect 319170 453218 319406 453454
rect 319170 452898 319406 453134
rect 349890 453218 350126 453454
rect 349890 452898 350126 453134
rect 380610 453218 380846 453454
rect 380610 452898 380846 453134
rect 411330 453218 411566 453454
rect 411330 452898 411566 453134
rect 442050 453218 442286 453454
rect 442050 452898 442286 453134
rect 472770 453218 473006 453454
rect 472770 452898 473006 453134
rect 503490 453218 503726 453454
rect 503490 452898 503726 453134
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 58050 435218 58286 435454
rect 58050 434898 58286 435134
rect 88770 435218 89006 435454
rect 88770 434898 89006 435134
rect 119490 435218 119726 435454
rect 119490 434898 119726 435134
rect 150210 435218 150446 435454
rect 150210 434898 150446 435134
rect 180930 435218 181166 435454
rect 180930 434898 181166 435134
rect 211650 435218 211886 435454
rect 211650 434898 211886 435134
rect 242370 435218 242606 435454
rect 242370 434898 242606 435134
rect 273090 435218 273326 435454
rect 273090 434898 273326 435134
rect 303810 435218 304046 435454
rect 303810 434898 304046 435134
rect 334530 435218 334766 435454
rect 334530 434898 334766 435134
rect 365250 435218 365486 435454
rect 365250 434898 365486 435134
rect 395970 435218 396206 435454
rect 395970 434898 396206 435134
rect 426690 435218 426926 435454
rect 426690 434898 426926 435134
rect 457410 435218 457646 435454
rect 457410 434898 457646 435134
rect 488130 435218 488366 435454
rect 488130 434898 488366 435134
rect 518850 435218 519086 435454
rect 518850 434898 519086 435134
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 73410 417218 73646 417454
rect 73410 416898 73646 417134
rect 104130 417218 104366 417454
rect 104130 416898 104366 417134
rect 134850 417218 135086 417454
rect 134850 416898 135086 417134
rect 165570 417218 165806 417454
rect 165570 416898 165806 417134
rect 196290 417218 196526 417454
rect 196290 416898 196526 417134
rect 227010 417218 227246 417454
rect 227010 416898 227246 417134
rect 257730 417218 257966 417454
rect 257730 416898 257966 417134
rect 288450 417218 288686 417454
rect 288450 416898 288686 417134
rect 319170 417218 319406 417454
rect 319170 416898 319406 417134
rect 349890 417218 350126 417454
rect 349890 416898 350126 417134
rect 380610 417218 380846 417454
rect 380610 416898 380846 417134
rect 411330 417218 411566 417454
rect 411330 416898 411566 417134
rect 442050 417218 442286 417454
rect 442050 416898 442286 417134
rect 472770 417218 473006 417454
rect 472770 416898 473006 417134
rect 503490 417218 503726 417454
rect 503490 416898 503726 417134
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 58050 399218 58286 399454
rect 58050 398898 58286 399134
rect 88770 399218 89006 399454
rect 88770 398898 89006 399134
rect 119490 399218 119726 399454
rect 119490 398898 119726 399134
rect 150210 399218 150446 399454
rect 150210 398898 150446 399134
rect 180930 399218 181166 399454
rect 180930 398898 181166 399134
rect 211650 399218 211886 399454
rect 211650 398898 211886 399134
rect 242370 399218 242606 399454
rect 242370 398898 242606 399134
rect 273090 399218 273326 399454
rect 273090 398898 273326 399134
rect 303810 399218 304046 399454
rect 303810 398898 304046 399134
rect 334530 399218 334766 399454
rect 334530 398898 334766 399134
rect 365250 399218 365486 399454
rect 365250 398898 365486 399134
rect 395970 399218 396206 399454
rect 395970 398898 396206 399134
rect 426690 399218 426926 399454
rect 426690 398898 426926 399134
rect 457410 399218 457646 399454
rect 457410 398898 457646 399134
rect 488130 399218 488366 399454
rect 488130 398898 488366 399134
rect 518850 399218 519086 399454
rect 518850 398898 519086 399134
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 73410 381218 73646 381454
rect 73410 380898 73646 381134
rect 104130 381218 104366 381454
rect 104130 380898 104366 381134
rect 134850 381218 135086 381454
rect 134850 380898 135086 381134
rect 165570 381218 165806 381454
rect 165570 380898 165806 381134
rect 196290 381218 196526 381454
rect 196290 380898 196526 381134
rect 227010 381218 227246 381454
rect 227010 380898 227246 381134
rect 257730 381218 257966 381454
rect 257730 380898 257966 381134
rect 288450 381218 288686 381454
rect 288450 380898 288686 381134
rect 319170 381218 319406 381454
rect 319170 380898 319406 381134
rect 349890 381218 350126 381454
rect 349890 380898 350126 381134
rect 380610 381218 380846 381454
rect 380610 380898 380846 381134
rect 411330 381218 411566 381454
rect 411330 380898 411566 381134
rect 442050 381218 442286 381454
rect 442050 380898 442286 381134
rect 472770 381218 473006 381454
rect 472770 380898 473006 381134
rect 503490 381218 503726 381454
rect 503490 380898 503726 381134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 58050 363218 58286 363454
rect 58050 362898 58286 363134
rect 88770 363218 89006 363454
rect 88770 362898 89006 363134
rect 119490 363218 119726 363454
rect 119490 362898 119726 363134
rect 150210 363218 150446 363454
rect 150210 362898 150446 363134
rect 180930 363218 181166 363454
rect 180930 362898 181166 363134
rect 211650 363218 211886 363454
rect 211650 362898 211886 363134
rect 242370 363218 242606 363454
rect 242370 362898 242606 363134
rect 273090 363218 273326 363454
rect 273090 362898 273326 363134
rect 303810 363218 304046 363454
rect 303810 362898 304046 363134
rect 334530 363218 334766 363454
rect 334530 362898 334766 363134
rect 365250 363218 365486 363454
rect 365250 362898 365486 363134
rect 395970 363218 396206 363454
rect 395970 362898 396206 363134
rect 426690 363218 426926 363454
rect 426690 362898 426926 363134
rect 457410 363218 457646 363454
rect 457410 362898 457646 363134
rect 488130 363218 488366 363454
rect 488130 362898 488366 363134
rect 518850 363218 519086 363454
rect 518850 362898 519086 363134
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 73410 345218 73646 345454
rect 73410 344898 73646 345134
rect 104130 345218 104366 345454
rect 104130 344898 104366 345134
rect 134850 345218 135086 345454
rect 134850 344898 135086 345134
rect 165570 345218 165806 345454
rect 165570 344898 165806 345134
rect 196290 345218 196526 345454
rect 196290 344898 196526 345134
rect 227010 345218 227246 345454
rect 227010 344898 227246 345134
rect 257730 345218 257966 345454
rect 257730 344898 257966 345134
rect 288450 345218 288686 345454
rect 288450 344898 288686 345134
rect 319170 345218 319406 345454
rect 319170 344898 319406 345134
rect 349890 345218 350126 345454
rect 349890 344898 350126 345134
rect 380610 345218 380846 345454
rect 380610 344898 380846 345134
rect 411330 345218 411566 345454
rect 411330 344898 411566 345134
rect 442050 345218 442286 345454
rect 442050 344898 442286 345134
rect 472770 345218 473006 345454
rect 472770 344898 473006 345134
rect 503490 345218 503726 345454
rect 503490 344898 503726 345134
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 58050 327218 58286 327454
rect 58050 326898 58286 327134
rect 88770 327218 89006 327454
rect 88770 326898 89006 327134
rect 119490 327218 119726 327454
rect 119490 326898 119726 327134
rect 150210 327218 150446 327454
rect 150210 326898 150446 327134
rect 180930 327218 181166 327454
rect 180930 326898 181166 327134
rect 211650 327218 211886 327454
rect 211650 326898 211886 327134
rect 242370 327218 242606 327454
rect 242370 326898 242606 327134
rect 273090 327218 273326 327454
rect 273090 326898 273326 327134
rect 303810 327218 304046 327454
rect 303810 326898 304046 327134
rect 334530 327218 334766 327454
rect 334530 326898 334766 327134
rect 365250 327218 365486 327454
rect 365250 326898 365486 327134
rect 395970 327218 396206 327454
rect 395970 326898 396206 327134
rect 426690 327218 426926 327454
rect 426690 326898 426926 327134
rect 457410 327218 457646 327454
rect 457410 326898 457646 327134
rect 488130 327218 488366 327454
rect 488130 326898 488366 327134
rect 518850 327218 519086 327454
rect 518850 326898 519086 327134
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 73410 309218 73646 309454
rect 73410 308898 73646 309134
rect 104130 309218 104366 309454
rect 104130 308898 104366 309134
rect 134850 309218 135086 309454
rect 134850 308898 135086 309134
rect 165570 309218 165806 309454
rect 165570 308898 165806 309134
rect 196290 309218 196526 309454
rect 196290 308898 196526 309134
rect 227010 309218 227246 309454
rect 227010 308898 227246 309134
rect 257730 309218 257966 309454
rect 257730 308898 257966 309134
rect 288450 309218 288686 309454
rect 288450 308898 288686 309134
rect 319170 309218 319406 309454
rect 319170 308898 319406 309134
rect 349890 309218 350126 309454
rect 349890 308898 350126 309134
rect 380610 309218 380846 309454
rect 380610 308898 380846 309134
rect 411330 309218 411566 309454
rect 411330 308898 411566 309134
rect 442050 309218 442286 309454
rect 442050 308898 442286 309134
rect 472770 309218 473006 309454
rect 472770 308898 473006 309134
rect 503490 309218 503726 309454
rect 503490 308898 503726 309134
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 58050 291218 58286 291454
rect 58050 290898 58286 291134
rect 88770 291218 89006 291454
rect 88770 290898 89006 291134
rect 119490 291218 119726 291454
rect 119490 290898 119726 291134
rect 150210 291218 150446 291454
rect 150210 290898 150446 291134
rect 180930 291218 181166 291454
rect 180930 290898 181166 291134
rect 211650 291218 211886 291454
rect 211650 290898 211886 291134
rect 242370 291218 242606 291454
rect 242370 290898 242606 291134
rect 273090 291218 273326 291454
rect 273090 290898 273326 291134
rect 303810 291218 304046 291454
rect 303810 290898 304046 291134
rect 334530 291218 334766 291454
rect 334530 290898 334766 291134
rect 365250 291218 365486 291454
rect 365250 290898 365486 291134
rect 395970 291218 396206 291454
rect 395970 290898 396206 291134
rect 426690 291218 426926 291454
rect 426690 290898 426926 291134
rect 457410 291218 457646 291454
rect 457410 290898 457646 291134
rect 488130 291218 488366 291454
rect 488130 290898 488366 291134
rect 518850 291218 519086 291454
rect 518850 290898 519086 291134
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 73410 273218 73646 273454
rect 73410 272898 73646 273134
rect 104130 273218 104366 273454
rect 104130 272898 104366 273134
rect 134850 273218 135086 273454
rect 134850 272898 135086 273134
rect 165570 273218 165806 273454
rect 165570 272898 165806 273134
rect 196290 273218 196526 273454
rect 196290 272898 196526 273134
rect 227010 273218 227246 273454
rect 227010 272898 227246 273134
rect 257730 273218 257966 273454
rect 257730 272898 257966 273134
rect 288450 273218 288686 273454
rect 288450 272898 288686 273134
rect 319170 273218 319406 273454
rect 319170 272898 319406 273134
rect 349890 273218 350126 273454
rect 349890 272898 350126 273134
rect 380610 273218 380846 273454
rect 380610 272898 380846 273134
rect 411330 273218 411566 273454
rect 411330 272898 411566 273134
rect 442050 273218 442286 273454
rect 442050 272898 442286 273134
rect 472770 273218 473006 273454
rect 472770 272898 473006 273134
rect 503490 273218 503726 273454
rect 503490 272898 503726 273134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 58050 255218 58286 255454
rect 58050 254898 58286 255134
rect 88770 255218 89006 255454
rect 88770 254898 89006 255134
rect 119490 255218 119726 255454
rect 119490 254898 119726 255134
rect 150210 255218 150446 255454
rect 150210 254898 150446 255134
rect 180930 255218 181166 255454
rect 180930 254898 181166 255134
rect 211650 255218 211886 255454
rect 211650 254898 211886 255134
rect 242370 255218 242606 255454
rect 242370 254898 242606 255134
rect 273090 255218 273326 255454
rect 273090 254898 273326 255134
rect 303810 255218 304046 255454
rect 303810 254898 304046 255134
rect 334530 255218 334766 255454
rect 334530 254898 334766 255134
rect 365250 255218 365486 255454
rect 365250 254898 365486 255134
rect 395970 255218 396206 255454
rect 395970 254898 396206 255134
rect 426690 255218 426926 255454
rect 426690 254898 426926 255134
rect 457410 255218 457646 255454
rect 457410 254898 457646 255134
rect 488130 255218 488366 255454
rect 488130 254898 488366 255134
rect 518850 255218 519086 255454
rect 518850 254898 519086 255134
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 73410 237218 73646 237454
rect 73410 236898 73646 237134
rect 104130 237218 104366 237454
rect 104130 236898 104366 237134
rect 134850 237218 135086 237454
rect 134850 236898 135086 237134
rect 165570 237218 165806 237454
rect 165570 236898 165806 237134
rect 196290 237218 196526 237454
rect 196290 236898 196526 237134
rect 227010 237218 227246 237454
rect 227010 236898 227246 237134
rect 257730 237218 257966 237454
rect 257730 236898 257966 237134
rect 288450 237218 288686 237454
rect 288450 236898 288686 237134
rect 319170 237218 319406 237454
rect 319170 236898 319406 237134
rect 349890 237218 350126 237454
rect 349890 236898 350126 237134
rect 380610 237218 380846 237454
rect 380610 236898 380846 237134
rect 411330 237218 411566 237454
rect 411330 236898 411566 237134
rect 442050 237218 442286 237454
rect 442050 236898 442286 237134
rect 472770 237218 473006 237454
rect 472770 236898 473006 237134
rect 503490 237218 503726 237454
rect 503490 236898 503726 237134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 58050 219218 58286 219454
rect 58050 218898 58286 219134
rect 88770 219218 89006 219454
rect 88770 218898 89006 219134
rect 119490 219218 119726 219454
rect 119490 218898 119726 219134
rect 150210 219218 150446 219454
rect 150210 218898 150446 219134
rect 180930 219218 181166 219454
rect 180930 218898 181166 219134
rect 211650 219218 211886 219454
rect 211650 218898 211886 219134
rect 242370 219218 242606 219454
rect 242370 218898 242606 219134
rect 273090 219218 273326 219454
rect 273090 218898 273326 219134
rect 303810 219218 304046 219454
rect 303810 218898 304046 219134
rect 334530 219218 334766 219454
rect 334530 218898 334766 219134
rect 365250 219218 365486 219454
rect 365250 218898 365486 219134
rect 395970 219218 396206 219454
rect 395970 218898 396206 219134
rect 426690 219218 426926 219454
rect 426690 218898 426926 219134
rect 457410 219218 457646 219454
rect 457410 218898 457646 219134
rect 488130 219218 488366 219454
rect 488130 218898 488366 219134
rect 518850 219218 519086 219454
rect 518850 218898 519086 219134
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 73410 201218 73646 201454
rect 73410 200898 73646 201134
rect 104130 201218 104366 201454
rect 104130 200898 104366 201134
rect 134850 201218 135086 201454
rect 134850 200898 135086 201134
rect 165570 201218 165806 201454
rect 165570 200898 165806 201134
rect 196290 201218 196526 201454
rect 196290 200898 196526 201134
rect 227010 201218 227246 201454
rect 227010 200898 227246 201134
rect 257730 201218 257966 201454
rect 257730 200898 257966 201134
rect 288450 201218 288686 201454
rect 288450 200898 288686 201134
rect 319170 201218 319406 201454
rect 319170 200898 319406 201134
rect 349890 201218 350126 201454
rect 349890 200898 350126 201134
rect 380610 201218 380846 201454
rect 380610 200898 380846 201134
rect 411330 201218 411566 201454
rect 411330 200898 411566 201134
rect 442050 201218 442286 201454
rect 442050 200898 442286 201134
rect 472770 201218 473006 201454
rect 472770 200898 473006 201134
rect 503490 201218 503726 201454
rect 503490 200898 503726 201134
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 58050 183218 58286 183454
rect 58050 182898 58286 183134
rect 88770 183218 89006 183454
rect 88770 182898 89006 183134
rect 119490 183218 119726 183454
rect 119490 182898 119726 183134
rect 150210 183218 150446 183454
rect 150210 182898 150446 183134
rect 180930 183218 181166 183454
rect 180930 182898 181166 183134
rect 211650 183218 211886 183454
rect 211650 182898 211886 183134
rect 242370 183218 242606 183454
rect 242370 182898 242606 183134
rect 273090 183218 273326 183454
rect 273090 182898 273326 183134
rect 303810 183218 304046 183454
rect 303810 182898 304046 183134
rect 334530 183218 334766 183454
rect 334530 182898 334766 183134
rect 365250 183218 365486 183454
rect 365250 182898 365486 183134
rect 395970 183218 396206 183454
rect 395970 182898 396206 183134
rect 426690 183218 426926 183454
rect 426690 182898 426926 183134
rect 457410 183218 457646 183454
rect 457410 182898 457646 183134
rect 488130 183218 488366 183454
rect 488130 182898 488366 183134
rect 518850 183218 519086 183454
rect 518850 182898 519086 183134
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 73410 165218 73646 165454
rect 73410 164898 73646 165134
rect 104130 165218 104366 165454
rect 104130 164898 104366 165134
rect 134850 165218 135086 165454
rect 134850 164898 135086 165134
rect 165570 165218 165806 165454
rect 165570 164898 165806 165134
rect 196290 165218 196526 165454
rect 196290 164898 196526 165134
rect 227010 165218 227246 165454
rect 227010 164898 227246 165134
rect 257730 165218 257966 165454
rect 257730 164898 257966 165134
rect 288450 165218 288686 165454
rect 288450 164898 288686 165134
rect 319170 165218 319406 165454
rect 319170 164898 319406 165134
rect 349890 165218 350126 165454
rect 349890 164898 350126 165134
rect 380610 165218 380846 165454
rect 380610 164898 380846 165134
rect 411330 165218 411566 165454
rect 411330 164898 411566 165134
rect 442050 165218 442286 165454
rect 442050 164898 442286 165134
rect 472770 165218 473006 165454
rect 472770 164898 473006 165134
rect 503490 165218 503726 165454
rect 503490 164898 503726 165134
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 58050 147218 58286 147454
rect 58050 146898 58286 147134
rect 88770 147218 89006 147454
rect 88770 146898 89006 147134
rect 119490 147218 119726 147454
rect 119490 146898 119726 147134
rect 150210 147218 150446 147454
rect 150210 146898 150446 147134
rect 180930 147218 181166 147454
rect 180930 146898 181166 147134
rect 211650 147218 211886 147454
rect 211650 146898 211886 147134
rect 242370 147218 242606 147454
rect 242370 146898 242606 147134
rect 273090 147218 273326 147454
rect 273090 146898 273326 147134
rect 303810 147218 304046 147454
rect 303810 146898 304046 147134
rect 334530 147218 334766 147454
rect 334530 146898 334766 147134
rect 365250 147218 365486 147454
rect 365250 146898 365486 147134
rect 395970 147218 396206 147454
rect 395970 146898 396206 147134
rect 426690 147218 426926 147454
rect 426690 146898 426926 147134
rect 457410 147218 457646 147454
rect 457410 146898 457646 147134
rect 488130 147218 488366 147454
rect 488130 146898 488366 147134
rect 518850 147218 519086 147454
rect 518850 146898 519086 147134
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 73410 129218 73646 129454
rect 73410 128898 73646 129134
rect 104130 129218 104366 129454
rect 104130 128898 104366 129134
rect 134850 129218 135086 129454
rect 134850 128898 135086 129134
rect 165570 129218 165806 129454
rect 165570 128898 165806 129134
rect 196290 129218 196526 129454
rect 196290 128898 196526 129134
rect 227010 129218 227246 129454
rect 227010 128898 227246 129134
rect 257730 129218 257966 129454
rect 257730 128898 257966 129134
rect 288450 129218 288686 129454
rect 288450 128898 288686 129134
rect 319170 129218 319406 129454
rect 319170 128898 319406 129134
rect 349890 129218 350126 129454
rect 349890 128898 350126 129134
rect 380610 129218 380846 129454
rect 380610 128898 380846 129134
rect 411330 129218 411566 129454
rect 411330 128898 411566 129134
rect 442050 129218 442286 129454
rect 442050 128898 442286 129134
rect 472770 129218 473006 129454
rect 472770 128898 473006 129134
rect 503490 129218 503726 129454
rect 503490 128898 503726 129134
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 58050 111218 58286 111454
rect 58050 110898 58286 111134
rect 88770 111218 89006 111454
rect 88770 110898 89006 111134
rect 119490 111218 119726 111454
rect 119490 110898 119726 111134
rect 150210 111218 150446 111454
rect 150210 110898 150446 111134
rect 180930 111218 181166 111454
rect 180930 110898 181166 111134
rect 211650 111218 211886 111454
rect 211650 110898 211886 111134
rect 242370 111218 242606 111454
rect 242370 110898 242606 111134
rect 273090 111218 273326 111454
rect 273090 110898 273326 111134
rect 303810 111218 304046 111454
rect 303810 110898 304046 111134
rect 334530 111218 334766 111454
rect 334530 110898 334766 111134
rect 365250 111218 365486 111454
rect 365250 110898 365486 111134
rect 395970 111218 396206 111454
rect 395970 110898 396206 111134
rect 426690 111218 426926 111454
rect 426690 110898 426926 111134
rect 457410 111218 457646 111454
rect 457410 110898 457646 111134
rect 488130 111218 488366 111454
rect 488130 110898 488366 111134
rect 518850 111218 519086 111454
rect 518850 110898 519086 111134
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 73410 93218 73646 93454
rect 73410 92898 73646 93134
rect 104130 93218 104366 93454
rect 104130 92898 104366 93134
rect 134850 93218 135086 93454
rect 134850 92898 135086 93134
rect 165570 93218 165806 93454
rect 165570 92898 165806 93134
rect 196290 93218 196526 93454
rect 196290 92898 196526 93134
rect 227010 93218 227246 93454
rect 227010 92898 227246 93134
rect 257730 93218 257966 93454
rect 257730 92898 257966 93134
rect 288450 93218 288686 93454
rect 288450 92898 288686 93134
rect 319170 93218 319406 93454
rect 319170 92898 319406 93134
rect 349890 93218 350126 93454
rect 349890 92898 350126 93134
rect 380610 93218 380846 93454
rect 380610 92898 380846 93134
rect 411330 93218 411566 93454
rect 411330 92898 411566 93134
rect 442050 93218 442286 93454
rect 442050 92898 442286 93134
rect 472770 93218 473006 93454
rect 472770 92898 473006 93134
rect 503490 93218 503726 93454
rect 503490 92898 503726 93134
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 58050 75218 58286 75454
rect 58050 74898 58286 75134
rect 88770 75218 89006 75454
rect 88770 74898 89006 75134
rect 119490 75218 119726 75454
rect 119490 74898 119726 75134
rect 150210 75218 150446 75454
rect 150210 74898 150446 75134
rect 180930 75218 181166 75454
rect 180930 74898 181166 75134
rect 211650 75218 211886 75454
rect 211650 74898 211886 75134
rect 242370 75218 242606 75454
rect 242370 74898 242606 75134
rect 273090 75218 273326 75454
rect 273090 74898 273326 75134
rect 303810 75218 304046 75454
rect 303810 74898 304046 75134
rect 334530 75218 334766 75454
rect 334530 74898 334766 75134
rect 365250 75218 365486 75454
rect 365250 74898 365486 75134
rect 395970 75218 396206 75454
rect 395970 74898 396206 75134
rect 426690 75218 426926 75454
rect 426690 74898 426926 75134
rect 457410 75218 457646 75454
rect 457410 74898 457646 75134
rect 488130 75218 488366 75454
rect 488130 74898 488366 75134
rect 518850 75218 519086 75454
rect 518850 74898 519086 75134
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 73410 633454
rect 73646 633218 104130 633454
rect 104366 633218 134850 633454
rect 135086 633218 165570 633454
rect 165806 633218 196290 633454
rect 196526 633218 227010 633454
rect 227246 633218 257730 633454
rect 257966 633218 288450 633454
rect 288686 633218 319170 633454
rect 319406 633218 349890 633454
rect 350126 633218 380610 633454
rect 380846 633218 411330 633454
rect 411566 633218 442050 633454
rect 442286 633218 472770 633454
rect 473006 633218 503490 633454
rect 503726 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 73410 633134
rect 73646 632898 104130 633134
rect 104366 632898 134850 633134
rect 135086 632898 165570 633134
rect 165806 632898 196290 633134
rect 196526 632898 227010 633134
rect 227246 632898 257730 633134
rect 257966 632898 288450 633134
rect 288686 632898 319170 633134
rect 319406 632898 349890 633134
rect 350126 632898 380610 633134
rect 380846 632898 411330 633134
rect 411566 632898 442050 633134
rect 442286 632898 472770 633134
rect 473006 632898 503490 633134
rect 503726 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 58050 615454
rect 58286 615218 88770 615454
rect 89006 615218 119490 615454
rect 119726 615218 150210 615454
rect 150446 615218 180930 615454
rect 181166 615218 211650 615454
rect 211886 615218 242370 615454
rect 242606 615218 273090 615454
rect 273326 615218 303810 615454
rect 304046 615218 334530 615454
rect 334766 615218 365250 615454
rect 365486 615218 395970 615454
rect 396206 615218 426690 615454
rect 426926 615218 457410 615454
rect 457646 615218 488130 615454
rect 488366 615218 518850 615454
rect 519086 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 58050 615134
rect 58286 614898 88770 615134
rect 89006 614898 119490 615134
rect 119726 614898 150210 615134
rect 150446 614898 180930 615134
rect 181166 614898 211650 615134
rect 211886 614898 242370 615134
rect 242606 614898 273090 615134
rect 273326 614898 303810 615134
rect 304046 614898 334530 615134
rect 334766 614898 365250 615134
rect 365486 614898 395970 615134
rect 396206 614898 426690 615134
rect 426926 614898 457410 615134
rect 457646 614898 488130 615134
rect 488366 614898 518850 615134
rect 519086 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 73410 597454
rect 73646 597218 104130 597454
rect 104366 597218 134850 597454
rect 135086 597218 165570 597454
rect 165806 597218 196290 597454
rect 196526 597218 227010 597454
rect 227246 597218 257730 597454
rect 257966 597218 288450 597454
rect 288686 597218 319170 597454
rect 319406 597218 349890 597454
rect 350126 597218 380610 597454
rect 380846 597218 411330 597454
rect 411566 597218 442050 597454
rect 442286 597218 472770 597454
rect 473006 597218 503490 597454
rect 503726 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 73410 597134
rect 73646 596898 104130 597134
rect 104366 596898 134850 597134
rect 135086 596898 165570 597134
rect 165806 596898 196290 597134
rect 196526 596898 227010 597134
rect 227246 596898 257730 597134
rect 257966 596898 288450 597134
rect 288686 596898 319170 597134
rect 319406 596898 349890 597134
rect 350126 596898 380610 597134
rect 380846 596898 411330 597134
rect 411566 596898 442050 597134
rect 442286 596898 472770 597134
rect 473006 596898 503490 597134
rect 503726 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 58050 579454
rect 58286 579218 88770 579454
rect 89006 579218 119490 579454
rect 119726 579218 150210 579454
rect 150446 579218 180930 579454
rect 181166 579218 211650 579454
rect 211886 579218 242370 579454
rect 242606 579218 273090 579454
rect 273326 579218 303810 579454
rect 304046 579218 334530 579454
rect 334766 579218 365250 579454
rect 365486 579218 395970 579454
rect 396206 579218 426690 579454
rect 426926 579218 457410 579454
rect 457646 579218 488130 579454
rect 488366 579218 518850 579454
rect 519086 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 58050 579134
rect 58286 578898 88770 579134
rect 89006 578898 119490 579134
rect 119726 578898 150210 579134
rect 150446 578898 180930 579134
rect 181166 578898 211650 579134
rect 211886 578898 242370 579134
rect 242606 578898 273090 579134
rect 273326 578898 303810 579134
rect 304046 578898 334530 579134
rect 334766 578898 365250 579134
rect 365486 578898 395970 579134
rect 396206 578898 426690 579134
rect 426926 578898 457410 579134
rect 457646 578898 488130 579134
rect 488366 578898 518850 579134
rect 519086 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 73410 561454
rect 73646 561218 104130 561454
rect 104366 561218 134850 561454
rect 135086 561218 165570 561454
rect 165806 561218 196290 561454
rect 196526 561218 227010 561454
rect 227246 561218 257730 561454
rect 257966 561218 288450 561454
rect 288686 561218 319170 561454
rect 319406 561218 349890 561454
rect 350126 561218 380610 561454
rect 380846 561218 411330 561454
rect 411566 561218 442050 561454
rect 442286 561218 472770 561454
rect 473006 561218 503490 561454
rect 503726 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 73410 561134
rect 73646 560898 104130 561134
rect 104366 560898 134850 561134
rect 135086 560898 165570 561134
rect 165806 560898 196290 561134
rect 196526 560898 227010 561134
rect 227246 560898 257730 561134
rect 257966 560898 288450 561134
rect 288686 560898 319170 561134
rect 319406 560898 349890 561134
rect 350126 560898 380610 561134
rect 380846 560898 411330 561134
rect 411566 560898 442050 561134
rect 442286 560898 472770 561134
rect 473006 560898 503490 561134
rect 503726 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 58050 543454
rect 58286 543218 88770 543454
rect 89006 543218 119490 543454
rect 119726 543218 150210 543454
rect 150446 543218 180930 543454
rect 181166 543218 211650 543454
rect 211886 543218 242370 543454
rect 242606 543218 273090 543454
rect 273326 543218 303810 543454
rect 304046 543218 334530 543454
rect 334766 543218 365250 543454
rect 365486 543218 395970 543454
rect 396206 543218 426690 543454
rect 426926 543218 457410 543454
rect 457646 543218 488130 543454
rect 488366 543218 518850 543454
rect 519086 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 58050 543134
rect 58286 542898 88770 543134
rect 89006 542898 119490 543134
rect 119726 542898 150210 543134
rect 150446 542898 180930 543134
rect 181166 542898 211650 543134
rect 211886 542898 242370 543134
rect 242606 542898 273090 543134
rect 273326 542898 303810 543134
rect 304046 542898 334530 543134
rect 334766 542898 365250 543134
rect 365486 542898 395970 543134
rect 396206 542898 426690 543134
rect 426926 542898 457410 543134
rect 457646 542898 488130 543134
rect 488366 542898 518850 543134
rect 519086 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 73410 525454
rect 73646 525218 104130 525454
rect 104366 525218 134850 525454
rect 135086 525218 165570 525454
rect 165806 525218 196290 525454
rect 196526 525218 227010 525454
rect 227246 525218 257730 525454
rect 257966 525218 288450 525454
rect 288686 525218 319170 525454
rect 319406 525218 349890 525454
rect 350126 525218 380610 525454
rect 380846 525218 411330 525454
rect 411566 525218 442050 525454
rect 442286 525218 472770 525454
rect 473006 525218 503490 525454
rect 503726 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 73410 525134
rect 73646 524898 104130 525134
rect 104366 524898 134850 525134
rect 135086 524898 165570 525134
rect 165806 524898 196290 525134
rect 196526 524898 227010 525134
rect 227246 524898 257730 525134
rect 257966 524898 288450 525134
rect 288686 524898 319170 525134
rect 319406 524898 349890 525134
rect 350126 524898 380610 525134
rect 380846 524898 411330 525134
rect 411566 524898 442050 525134
rect 442286 524898 472770 525134
rect 473006 524898 503490 525134
rect 503726 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 58050 507454
rect 58286 507218 88770 507454
rect 89006 507218 119490 507454
rect 119726 507218 150210 507454
rect 150446 507218 180930 507454
rect 181166 507218 211650 507454
rect 211886 507218 242370 507454
rect 242606 507218 273090 507454
rect 273326 507218 303810 507454
rect 304046 507218 334530 507454
rect 334766 507218 365250 507454
rect 365486 507218 395970 507454
rect 396206 507218 426690 507454
rect 426926 507218 457410 507454
rect 457646 507218 488130 507454
rect 488366 507218 518850 507454
rect 519086 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 58050 507134
rect 58286 506898 88770 507134
rect 89006 506898 119490 507134
rect 119726 506898 150210 507134
rect 150446 506898 180930 507134
rect 181166 506898 211650 507134
rect 211886 506898 242370 507134
rect 242606 506898 273090 507134
rect 273326 506898 303810 507134
rect 304046 506898 334530 507134
rect 334766 506898 365250 507134
rect 365486 506898 395970 507134
rect 396206 506898 426690 507134
rect 426926 506898 457410 507134
rect 457646 506898 488130 507134
rect 488366 506898 518850 507134
rect 519086 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 73410 489454
rect 73646 489218 104130 489454
rect 104366 489218 134850 489454
rect 135086 489218 165570 489454
rect 165806 489218 196290 489454
rect 196526 489218 227010 489454
rect 227246 489218 257730 489454
rect 257966 489218 288450 489454
rect 288686 489218 319170 489454
rect 319406 489218 349890 489454
rect 350126 489218 380610 489454
rect 380846 489218 411330 489454
rect 411566 489218 442050 489454
rect 442286 489218 472770 489454
rect 473006 489218 503490 489454
rect 503726 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 73410 489134
rect 73646 488898 104130 489134
rect 104366 488898 134850 489134
rect 135086 488898 165570 489134
rect 165806 488898 196290 489134
rect 196526 488898 227010 489134
rect 227246 488898 257730 489134
rect 257966 488898 288450 489134
rect 288686 488898 319170 489134
rect 319406 488898 349890 489134
rect 350126 488898 380610 489134
rect 380846 488898 411330 489134
rect 411566 488898 442050 489134
rect 442286 488898 472770 489134
rect 473006 488898 503490 489134
rect 503726 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 58050 471454
rect 58286 471218 88770 471454
rect 89006 471218 119490 471454
rect 119726 471218 150210 471454
rect 150446 471218 180930 471454
rect 181166 471218 211650 471454
rect 211886 471218 242370 471454
rect 242606 471218 273090 471454
rect 273326 471218 303810 471454
rect 304046 471218 334530 471454
rect 334766 471218 365250 471454
rect 365486 471218 395970 471454
rect 396206 471218 426690 471454
rect 426926 471218 457410 471454
rect 457646 471218 488130 471454
rect 488366 471218 518850 471454
rect 519086 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 58050 471134
rect 58286 470898 88770 471134
rect 89006 470898 119490 471134
rect 119726 470898 150210 471134
rect 150446 470898 180930 471134
rect 181166 470898 211650 471134
rect 211886 470898 242370 471134
rect 242606 470898 273090 471134
rect 273326 470898 303810 471134
rect 304046 470898 334530 471134
rect 334766 470898 365250 471134
rect 365486 470898 395970 471134
rect 396206 470898 426690 471134
rect 426926 470898 457410 471134
rect 457646 470898 488130 471134
rect 488366 470898 518850 471134
rect 519086 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 73410 453454
rect 73646 453218 104130 453454
rect 104366 453218 134850 453454
rect 135086 453218 165570 453454
rect 165806 453218 196290 453454
rect 196526 453218 227010 453454
rect 227246 453218 257730 453454
rect 257966 453218 288450 453454
rect 288686 453218 319170 453454
rect 319406 453218 349890 453454
rect 350126 453218 380610 453454
rect 380846 453218 411330 453454
rect 411566 453218 442050 453454
rect 442286 453218 472770 453454
rect 473006 453218 503490 453454
rect 503726 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 73410 453134
rect 73646 452898 104130 453134
rect 104366 452898 134850 453134
rect 135086 452898 165570 453134
rect 165806 452898 196290 453134
rect 196526 452898 227010 453134
rect 227246 452898 257730 453134
rect 257966 452898 288450 453134
rect 288686 452898 319170 453134
rect 319406 452898 349890 453134
rect 350126 452898 380610 453134
rect 380846 452898 411330 453134
rect 411566 452898 442050 453134
rect 442286 452898 472770 453134
rect 473006 452898 503490 453134
rect 503726 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 58050 435454
rect 58286 435218 88770 435454
rect 89006 435218 119490 435454
rect 119726 435218 150210 435454
rect 150446 435218 180930 435454
rect 181166 435218 211650 435454
rect 211886 435218 242370 435454
rect 242606 435218 273090 435454
rect 273326 435218 303810 435454
rect 304046 435218 334530 435454
rect 334766 435218 365250 435454
rect 365486 435218 395970 435454
rect 396206 435218 426690 435454
rect 426926 435218 457410 435454
rect 457646 435218 488130 435454
rect 488366 435218 518850 435454
rect 519086 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 58050 435134
rect 58286 434898 88770 435134
rect 89006 434898 119490 435134
rect 119726 434898 150210 435134
rect 150446 434898 180930 435134
rect 181166 434898 211650 435134
rect 211886 434898 242370 435134
rect 242606 434898 273090 435134
rect 273326 434898 303810 435134
rect 304046 434898 334530 435134
rect 334766 434898 365250 435134
rect 365486 434898 395970 435134
rect 396206 434898 426690 435134
rect 426926 434898 457410 435134
rect 457646 434898 488130 435134
rect 488366 434898 518850 435134
rect 519086 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 73410 417454
rect 73646 417218 104130 417454
rect 104366 417218 134850 417454
rect 135086 417218 165570 417454
rect 165806 417218 196290 417454
rect 196526 417218 227010 417454
rect 227246 417218 257730 417454
rect 257966 417218 288450 417454
rect 288686 417218 319170 417454
rect 319406 417218 349890 417454
rect 350126 417218 380610 417454
rect 380846 417218 411330 417454
rect 411566 417218 442050 417454
rect 442286 417218 472770 417454
rect 473006 417218 503490 417454
rect 503726 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 73410 417134
rect 73646 416898 104130 417134
rect 104366 416898 134850 417134
rect 135086 416898 165570 417134
rect 165806 416898 196290 417134
rect 196526 416898 227010 417134
rect 227246 416898 257730 417134
rect 257966 416898 288450 417134
rect 288686 416898 319170 417134
rect 319406 416898 349890 417134
rect 350126 416898 380610 417134
rect 380846 416898 411330 417134
rect 411566 416898 442050 417134
rect 442286 416898 472770 417134
rect 473006 416898 503490 417134
rect 503726 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 58050 399454
rect 58286 399218 88770 399454
rect 89006 399218 119490 399454
rect 119726 399218 150210 399454
rect 150446 399218 180930 399454
rect 181166 399218 211650 399454
rect 211886 399218 242370 399454
rect 242606 399218 273090 399454
rect 273326 399218 303810 399454
rect 304046 399218 334530 399454
rect 334766 399218 365250 399454
rect 365486 399218 395970 399454
rect 396206 399218 426690 399454
rect 426926 399218 457410 399454
rect 457646 399218 488130 399454
rect 488366 399218 518850 399454
rect 519086 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 58050 399134
rect 58286 398898 88770 399134
rect 89006 398898 119490 399134
rect 119726 398898 150210 399134
rect 150446 398898 180930 399134
rect 181166 398898 211650 399134
rect 211886 398898 242370 399134
rect 242606 398898 273090 399134
rect 273326 398898 303810 399134
rect 304046 398898 334530 399134
rect 334766 398898 365250 399134
rect 365486 398898 395970 399134
rect 396206 398898 426690 399134
rect 426926 398898 457410 399134
rect 457646 398898 488130 399134
rect 488366 398898 518850 399134
rect 519086 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 73410 381454
rect 73646 381218 104130 381454
rect 104366 381218 134850 381454
rect 135086 381218 165570 381454
rect 165806 381218 196290 381454
rect 196526 381218 227010 381454
rect 227246 381218 257730 381454
rect 257966 381218 288450 381454
rect 288686 381218 319170 381454
rect 319406 381218 349890 381454
rect 350126 381218 380610 381454
rect 380846 381218 411330 381454
rect 411566 381218 442050 381454
rect 442286 381218 472770 381454
rect 473006 381218 503490 381454
rect 503726 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 73410 381134
rect 73646 380898 104130 381134
rect 104366 380898 134850 381134
rect 135086 380898 165570 381134
rect 165806 380898 196290 381134
rect 196526 380898 227010 381134
rect 227246 380898 257730 381134
rect 257966 380898 288450 381134
rect 288686 380898 319170 381134
rect 319406 380898 349890 381134
rect 350126 380898 380610 381134
rect 380846 380898 411330 381134
rect 411566 380898 442050 381134
rect 442286 380898 472770 381134
rect 473006 380898 503490 381134
rect 503726 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 58050 363454
rect 58286 363218 88770 363454
rect 89006 363218 119490 363454
rect 119726 363218 150210 363454
rect 150446 363218 180930 363454
rect 181166 363218 211650 363454
rect 211886 363218 242370 363454
rect 242606 363218 273090 363454
rect 273326 363218 303810 363454
rect 304046 363218 334530 363454
rect 334766 363218 365250 363454
rect 365486 363218 395970 363454
rect 396206 363218 426690 363454
rect 426926 363218 457410 363454
rect 457646 363218 488130 363454
rect 488366 363218 518850 363454
rect 519086 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 58050 363134
rect 58286 362898 88770 363134
rect 89006 362898 119490 363134
rect 119726 362898 150210 363134
rect 150446 362898 180930 363134
rect 181166 362898 211650 363134
rect 211886 362898 242370 363134
rect 242606 362898 273090 363134
rect 273326 362898 303810 363134
rect 304046 362898 334530 363134
rect 334766 362898 365250 363134
rect 365486 362898 395970 363134
rect 396206 362898 426690 363134
rect 426926 362898 457410 363134
rect 457646 362898 488130 363134
rect 488366 362898 518850 363134
rect 519086 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 73410 345454
rect 73646 345218 104130 345454
rect 104366 345218 134850 345454
rect 135086 345218 165570 345454
rect 165806 345218 196290 345454
rect 196526 345218 227010 345454
rect 227246 345218 257730 345454
rect 257966 345218 288450 345454
rect 288686 345218 319170 345454
rect 319406 345218 349890 345454
rect 350126 345218 380610 345454
rect 380846 345218 411330 345454
rect 411566 345218 442050 345454
rect 442286 345218 472770 345454
rect 473006 345218 503490 345454
rect 503726 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 73410 345134
rect 73646 344898 104130 345134
rect 104366 344898 134850 345134
rect 135086 344898 165570 345134
rect 165806 344898 196290 345134
rect 196526 344898 227010 345134
rect 227246 344898 257730 345134
rect 257966 344898 288450 345134
rect 288686 344898 319170 345134
rect 319406 344898 349890 345134
rect 350126 344898 380610 345134
rect 380846 344898 411330 345134
rect 411566 344898 442050 345134
rect 442286 344898 472770 345134
rect 473006 344898 503490 345134
rect 503726 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 58050 327454
rect 58286 327218 88770 327454
rect 89006 327218 119490 327454
rect 119726 327218 150210 327454
rect 150446 327218 180930 327454
rect 181166 327218 211650 327454
rect 211886 327218 242370 327454
rect 242606 327218 273090 327454
rect 273326 327218 303810 327454
rect 304046 327218 334530 327454
rect 334766 327218 365250 327454
rect 365486 327218 395970 327454
rect 396206 327218 426690 327454
rect 426926 327218 457410 327454
rect 457646 327218 488130 327454
rect 488366 327218 518850 327454
rect 519086 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 58050 327134
rect 58286 326898 88770 327134
rect 89006 326898 119490 327134
rect 119726 326898 150210 327134
rect 150446 326898 180930 327134
rect 181166 326898 211650 327134
rect 211886 326898 242370 327134
rect 242606 326898 273090 327134
rect 273326 326898 303810 327134
rect 304046 326898 334530 327134
rect 334766 326898 365250 327134
rect 365486 326898 395970 327134
rect 396206 326898 426690 327134
rect 426926 326898 457410 327134
rect 457646 326898 488130 327134
rect 488366 326898 518850 327134
rect 519086 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 73410 309454
rect 73646 309218 104130 309454
rect 104366 309218 134850 309454
rect 135086 309218 165570 309454
rect 165806 309218 196290 309454
rect 196526 309218 227010 309454
rect 227246 309218 257730 309454
rect 257966 309218 288450 309454
rect 288686 309218 319170 309454
rect 319406 309218 349890 309454
rect 350126 309218 380610 309454
rect 380846 309218 411330 309454
rect 411566 309218 442050 309454
rect 442286 309218 472770 309454
rect 473006 309218 503490 309454
rect 503726 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 73410 309134
rect 73646 308898 104130 309134
rect 104366 308898 134850 309134
rect 135086 308898 165570 309134
rect 165806 308898 196290 309134
rect 196526 308898 227010 309134
rect 227246 308898 257730 309134
rect 257966 308898 288450 309134
rect 288686 308898 319170 309134
rect 319406 308898 349890 309134
rect 350126 308898 380610 309134
rect 380846 308898 411330 309134
rect 411566 308898 442050 309134
rect 442286 308898 472770 309134
rect 473006 308898 503490 309134
rect 503726 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 58050 291454
rect 58286 291218 88770 291454
rect 89006 291218 119490 291454
rect 119726 291218 150210 291454
rect 150446 291218 180930 291454
rect 181166 291218 211650 291454
rect 211886 291218 242370 291454
rect 242606 291218 273090 291454
rect 273326 291218 303810 291454
rect 304046 291218 334530 291454
rect 334766 291218 365250 291454
rect 365486 291218 395970 291454
rect 396206 291218 426690 291454
rect 426926 291218 457410 291454
rect 457646 291218 488130 291454
rect 488366 291218 518850 291454
rect 519086 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 58050 291134
rect 58286 290898 88770 291134
rect 89006 290898 119490 291134
rect 119726 290898 150210 291134
rect 150446 290898 180930 291134
rect 181166 290898 211650 291134
rect 211886 290898 242370 291134
rect 242606 290898 273090 291134
rect 273326 290898 303810 291134
rect 304046 290898 334530 291134
rect 334766 290898 365250 291134
rect 365486 290898 395970 291134
rect 396206 290898 426690 291134
rect 426926 290898 457410 291134
rect 457646 290898 488130 291134
rect 488366 290898 518850 291134
rect 519086 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 73410 273454
rect 73646 273218 104130 273454
rect 104366 273218 134850 273454
rect 135086 273218 165570 273454
rect 165806 273218 196290 273454
rect 196526 273218 227010 273454
rect 227246 273218 257730 273454
rect 257966 273218 288450 273454
rect 288686 273218 319170 273454
rect 319406 273218 349890 273454
rect 350126 273218 380610 273454
rect 380846 273218 411330 273454
rect 411566 273218 442050 273454
rect 442286 273218 472770 273454
rect 473006 273218 503490 273454
rect 503726 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 73410 273134
rect 73646 272898 104130 273134
rect 104366 272898 134850 273134
rect 135086 272898 165570 273134
rect 165806 272898 196290 273134
rect 196526 272898 227010 273134
rect 227246 272898 257730 273134
rect 257966 272898 288450 273134
rect 288686 272898 319170 273134
rect 319406 272898 349890 273134
rect 350126 272898 380610 273134
rect 380846 272898 411330 273134
rect 411566 272898 442050 273134
rect 442286 272898 472770 273134
rect 473006 272898 503490 273134
rect 503726 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 58050 255454
rect 58286 255218 88770 255454
rect 89006 255218 119490 255454
rect 119726 255218 150210 255454
rect 150446 255218 180930 255454
rect 181166 255218 211650 255454
rect 211886 255218 242370 255454
rect 242606 255218 273090 255454
rect 273326 255218 303810 255454
rect 304046 255218 334530 255454
rect 334766 255218 365250 255454
rect 365486 255218 395970 255454
rect 396206 255218 426690 255454
rect 426926 255218 457410 255454
rect 457646 255218 488130 255454
rect 488366 255218 518850 255454
rect 519086 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 58050 255134
rect 58286 254898 88770 255134
rect 89006 254898 119490 255134
rect 119726 254898 150210 255134
rect 150446 254898 180930 255134
rect 181166 254898 211650 255134
rect 211886 254898 242370 255134
rect 242606 254898 273090 255134
rect 273326 254898 303810 255134
rect 304046 254898 334530 255134
rect 334766 254898 365250 255134
rect 365486 254898 395970 255134
rect 396206 254898 426690 255134
rect 426926 254898 457410 255134
rect 457646 254898 488130 255134
rect 488366 254898 518850 255134
rect 519086 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 73410 237454
rect 73646 237218 104130 237454
rect 104366 237218 134850 237454
rect 135086 237218 165570 237454
rect 165806 237218 196290 237454
rect 196526 237218 227010 237454
rect 227246 237218 257730 237454
rect 257966 237218 288450 237454
rect 288686 237218 319170 237454
rect 319406 237218 349890 237454
rect 350126 237218 380610 237454
rect 380846 237218 411330 237454
rect 411566 237218 442050 237454
rect 442286 237218 472770 237454
rect 473006 237218 503490 237454
rect 503726 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 73410 237134
rect 73646 236898 104130 237134
rect 104366 236898 134850 237134
rect 135086 236898 165570 237134
rect 165806 236898 196290 237134
rect 196526 236898 227010 237134
rect 227246 236898 257730 237134
rect 257966 236898 288450 237134
rect 288686 236898 319170 237134
rect 319406 236898 349890 237134
rect 350126 236898 380610 237134
rect 380846 236898 411330 237134
rect 411566 236898 442050 237134
rect 442286 236898 472770 237134
rect 473006 236898 503490 237134
rect 503726 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 58050 219454
rect 58286 219218 88770 219454
rect 89006 219218 119490 219454
rect 119726 219218 150210 219454
rect 150446 219218 180930 219454
rect 181166 219218 211650 219454
rect 211886 219218 242370 219454
rect 242606 219218 273090 219454
rect 273326 219218 303810 219454
rect 304046 219218 334530 219454
rect 334766 219218 365250 219454
rect 365486 219218 395970 219454
rect 396206 219218 426690 219454
rect 426926 219218 457410 219454
rect 457646 219218 488130 219454
rect 488366 219218 518850 219454
rect 519086 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 58050 219134
rect 58286 218898 88770 219134
rect 89006 218898 119490 219134
rect 119726 218898 150210 219134
rect 150446 218898 180930 219134
rect 181166 218898 211650 219134
rect 211886 218898 242370 219134
rect 242606 218898 273090 219134
rect 273326 218898 303810 219134
rect 304046 218898 334530 219134
rect 334766 218898 365250 219134
rect 365486 218898 395970 219134
rect 396206 218898 426690 219134
rect 426926 218898 457410 219134
rect 457646 218898 488130 219134
rect 488366 218898 518850 219134
rect 519086 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 73410 201454
rect 73646 201218 104130 201454
rect 104366 201218 134850 201454
rect 135086 201218 165570 201454
rect 165806 201218 196290 201454
rect 196526 201218 227010 201454
rect 227246 201218 257730 201454
rect 257966 201218 288450 201454
rect 288686 201218 319170 201454
rect 319406 201218 349890 201454
rect 350126 201218 380610 201454
rect 380846 201218 411330 201454
rect 411566 201218 442050 201454
rect 442286 201218 472770 201454
rect 473006 201218 503490 201454
rect 503726 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 73410 201134
rect 73646 200898 104130 201134
rect 104366 200898 134850 201134
rect 135086 200898 165570 201134
rect 165806 200898 196290 201134
rect 196526 200898 227010 201134
rect 227246 200898 257730 201134
rect 257966 200898 288450 201134
rect 288686 200898 319170 201134
rect 319406 200898 349890 201134
rect 350126 200898 380610 201134
rect 380846 200898 411330 201134
rect 411566 200898 442050 201134
rect 442286 200898 472770 201134
rect 473006 200898 503490 201134
rect 503726 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 58050 183454
rect 58286 183218 88770 183454
rect 89006 183218 119490 183454
rect 119726 183218 150210 183454
rect 150446 183218 180930 183454
rect 181166 183218 211650 183454
rect 211886 183218 242370 183454
rect 242606 183218 273090 183454
rect 273326 183218 303810 183454
rect 304046 183218 334530 183454
rect 334766 183218 365250 183454
rect 365486 183218 395970 183454
rect 396206 183218 426690 183454
rect 426926 183218 457410 183454
rect 457646 183218 488130 183454
rect 488366 183218 518850 183454
rect 519086 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 58050 183134
rect 58286 182898 88770 183134
rect 89006 182898 119490 183134
rect 119726 182898 150210 183134
rect 150446 182898 180930 183134
rect 181166 182898 211650 183134
rect 211886 182898 242370 183134
rect 242606 182898 273090 183134
rect 273326 182898 303810 183134
rect 304046 182898 334530 183134
rect 334766 182898 365250 183134
rect 365486 182898 395970 183134
rect 396206 182898 426690 183134
rect 426926 182898 457410 183134
rect 457646 182898 488130 183134
rect 488366 182898 518850 183134
rect 519086 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 73410 165454
rect 73646 165218 104130 165454
rect 104366 165218 134850 165454
rect 135086 165218 165570 165454
rect 165806 165218 196290 165454
rect 196526 165218 227010 165454
rect 227246 165218 257730 165454
rect 257966 165218 288450 165454
rect 288686 165218 319170 165454
rect 319406 165218 349890 165454
rect 350126 165218 380610 165454
rect 380846 165218 411330 165454
rect 411566 165218 442050 165454
rect 442286 165218 472770 165454
rect 473006 165218 503490 165454
rect 503726 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 73410 165134
rect 73646 164898 104130 165134
rect 104366 164898 134850 165134
rect 135086 164898 165570 165134
rect 165806 164898 196290 165134
rect 196526 164898 227010 165134
rect 227246 164898 257730 165134
rect 257966 164898 288450 165134
rect 288686 164898 319170 165134
rect 319406 164898 349890 165134
rect 350126 164898 380610 165134
rect 380846 164898 411330 165134
rect 411566 164898 442050 165134
rect 442286 164898 472770 165134
rect 473006 164898 503490 165134
rect 503726 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 58050 147454
rect 58286 147218 88770 147454
rect 89006 147218 119490 147454
rect 119726 147218 150210 147454
rect 150446 147218 180930 147454
rect 181166 147218 211650 147454
rect 211886 147218 242370 147454
rect 242606 147218 273090 147454
rect 273326 147218 303810 147454
rect 304046 147218 334530 147454
rect 334766 147218 365250 147454
rect 365486 147218 395970 147454
rect 396206 147218 426690 147454
rect 426926 147218 457410 147454
rect 457646 147218 488130 147454
rect 488366 147218 518850 147454
rect 519086 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 58050 147134
rect 58286 146898 88770 147134
rect 89006 146898 119490 147134
rect 119726 146898 150210 147134
rect 150446 146898 180930 147134
rect 181166 146898 211650 147134
rect 211886 146898 242370 147134
rect 242606 146898 273090 147134
rect 273326 146898 303810 147134
rect 304046 146898 334530 147134
rect 334766 146898 365250 147134
rect 365486 146898 395970 147134
rect 396206 146898 426690 147134
rect 426926 146898 457410 147134
rect 457646 146898 488130 147134
rect 488366 146898 518850 147134
rect 519086 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 73410 129454
rect 73646 129218 104130 129454
rect 104366 129218 134850 129454
rect 135086 129218 165570 129454
rect 165806 129218 196290 129454
rect 196526 129218 227010 129454
rect 227246 129218 257730 129454
rect 257966 129218 288450 129454
rect 288686 129218 319170 129454
rect 319406 129218 349890 129454
rect 350126 129218 380610 129454
rect 380846 129218 411330 129454
rect 411566 129218 442050 129454
rect 442286 129218 472770 129454
rect 473006 129218 503490 129454
rect 503726 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 73410 129134
rect 73646 128898 104130 129134
rect 104366 128898 134850 129134
rect 135086 128898 165570 129134
rect 165806 128898 196290 129134
rect 196526 128898 227010 129134
rect 227246 128898 257730 129134
rect 257966 128898 288450 129134
rect 288686 128898 319170 129134
rect 319406 128898 349890 129134
rect 350126 128898 380610 129134
rect 380846 128898 411330 129134
rect 411566 128898 442050 129134
rect 442286 128898 472770 129134
rect 473006 128898 503490 129134
rect 503726 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 58050 111454
rect 58286 111218 88770 111454
rect 89006 111218 119490 111454
rect 119726 111218 150210 111454
rect 150446 111218 180930 111454
rect 181166 111218 211650 111454
rect 211886 111218 242370 111454
rect 242606 111218 273090 111454
rect 273326 111218 303810 111454
rect 304046 111218 334530 111454
rect 334766 111218 365250 111454
rect 365486 111218 395970 111454
rect 396206 111218 426690 111454
rect 426926 111218 457410 111454
rect 457646 111218 488130 111454
rect 488366 111218 518850 111454
rect 519086 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 58050 111134
rect 58286 110898 88770 111134
rect 89006 110898 119490 111134
rect 119726 110898 150210 111134
rect 150446 110898 180930 111134
rect 181166 110898 211650 111134
rect 211886 110898 242370 111134
rect 242606 110898 273090 111134
rect 273326 110898 303810 111134
rect 304046 110898 334530 111134
rect 334766 110898 365250 111134
rect 365486 110898 395970 111134
rect 396206 110898 426690 111134
rect 426926 110898 457410 111134
rect 457646 110898 488130 111134
rect 488366 110898 518850 111134
rect 519086 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 73410 93454
rect 73646 93218 104130 93454
rect 104366 93218 134850 93454
rect 135086 93218 165570 93454
rect 165806 93218 196290 93454
rect 196526 93218 227010 93454
rect 227246 93218 257730 93454
rect 257966 93218 288450 93454
rect 288686 93218 319170 93454
rect 319406 93218 349890 93454
rect 350126 93218 380610 93454
rect 380846 93218 411330 93454
rect 411566 93218 442050 93454
rect 442286 93218 472770 93454
rect 473006 93218 503490 93454
rect 503726 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 73410 93134
rect 73646 92898 104130 93134
rect 104366 92898 134850 93134
rect 135086 92898 165570 93134
rect 165806 92898 196290 93134
rect 196526 92898 227010 93134
rect 227246 92898 257730 93134
rect 257966 92898 288450 93134
rect 288686 92898 319170 93134
rect 319406 92898 349890 93134
rect 350126 92898 380610 93134
rect 380846 92898 411330 93134
rect 411566 92898 442050 93134
rect 442286 92898 472770 93134
rect 473006 92898 503490 93134
rect 503726 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 58050 75454
rect 58286 75218 88770 75454
rect 89006 75218 119490 75454
rect 119726 75218 150210 75454
rect 150446 75218 180930 75454
rect 181166 75218 211650 75454
rect 211886 75218 242370 75454
rect 242606 75218 273090 75454
rect 273326 75218 303810 75454
rect 304046 75218 334530 75454
rect 334766 75218 365250 75454
rect 365486 75218 395970 75454
rect 396206 75218 426690 75454
rect 426926 75218 457410 75454
rect 457646 75218 488130 75454
rect 488366 75218 518850 75454
rect 519086 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 58050 75134
rect 58286 74898 88770 75134
rect 89006 74898 119490 75134
rect 119726 74898 150210 75134
rect 150446 74898 180930 75134
rect 181166 74898 211650 75134
rect 211886 74898 242370 75134
rect 242606 74898 273090 75134
rect 273326 74898 303810 75134
rect 304046 74898 334530 75134
rect 334766 74898 365250 75134
rect 365486 74898 395970 75134
rect 396206 74898 426690 75134
rect 426926 74898 457410 75134
rect 457646 74898 488130 75134
rect 488366 74898 518850 75134
rect 519086 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1636885634
transform 1 0 53800 0 1 65400
box 474 0 475899 573151
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 63400 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 640551 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 640551 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 640551 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 640551 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 640551 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 640551 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 640551 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 640551 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 640551 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 640551 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 640551 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 640551 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 640551 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 63400 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 640551 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 640551 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 640551 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 640551 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 640551 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 640551 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 640551 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 640551 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 640551 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 640551 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 640551 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 640551 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 640551 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 63400 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 640551 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 640551 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 640551 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 640551 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 640551 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 640551 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 640551 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 640551 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 640551 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 640551 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 640551 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 640551 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 640551 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 63400 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 640551 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 640551 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 640551 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 640551 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 640551 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 640551 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 640551 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 640551 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 640551 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 640551 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 640551 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 640551 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 640551 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 63400 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 640551 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 640551 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 640551 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 640551 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 640551 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 640551 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 640551 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 640551 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 640551 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 640551 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 640551 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 640551 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 640551 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 640551 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 63400 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 640551 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 640551 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 640551 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 640551 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 640551 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 640551 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 640551 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 640551 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 640551 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 640551 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 640551 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 640551 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 640551 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 63400 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 640551 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 640551 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 640551 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 640551 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 640551 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 640551 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 640551 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 640551 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 640551 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 640551 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 640551 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 640551 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 640551 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 640551 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 63400 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 640551 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 640551 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 640551 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 640551 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 640551 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 640551 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 640551 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 640551 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 640551 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 640551 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 640551 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 640551 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 640551 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 640551 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
