magic
tech sky130A
magscale 1 2
timestamp 1636880886
<< obsli1 >>
rect 1104 1309 475887 570673
<< obsm1 >>
rect 474 8 475899 570704
<< metal2 >>
rect 2042 572351 2098 573151
rect 6182 572351 6238 573151
rect 10322 572351 10378 573151
rect 14554 572351 14610 573151
rect 18694 572351 18750 573151
rect 22926 572351 22982 573151
rect 27066 572351 27122 573151
rect 31206 572351 31262 573151
rect 35438 572351 35494 573151
rect 39578 572351 39634 573151
rect 43810 572351 43866 573151
rect 47950 572351 48006 573151
rect 52090 572351 52146 573151
rect 56322 572351 56378 573151
rect 60462 572351 60518 573151
rect 64694 572351 64750 573151
rect 68834 572351 68890 573151
rect 72974 572351 73030 573151
rect 77206 572351 77262 573151
rect 81346 572351 81402 573151
rect 85578 572351 85634 573151
rect 89718 572351 89774 573151
rect 93858 572351 93914 573151
rect 98090 572351 98146 573151
rect 102230 572351 102286 573151
rect 106462 572351 106518 573151
rect 110602 572351 110658 573151
rect 114742 572351 114798 573151
rect 118974 572351 119030 573151
rect 123114 572351 123170 573151
rect 127346 572351 127402 573151
rect 131486 572351 131542 573151
rect 135626 572351 135682 573151
rect 139858 572351 139914 573151
rect 143998 572351 144054 573151
rect 148230 572351 148286 573151
rect 152370 572351 152426 573151
rect 156510 572351 156566 573151
rect 160742 572351 160798 573151
rect 164882 572351 164938 573151
rect 169114 572351 169170 573151
rect 173254 572351 173310 573151
rect 177394 572351 177450 573151
rect 181626 572351 181682 573151
rect 185766 572351 185822 573151
rect 189998 572351 190054 573151
rect 194138 572351 194194 573151
rect 198278 572351 198334 573151
rect 202510 572351 202566 573151
rect 206650 572351 206706 573151
rect 210882 572351 210938 573151
rect 215022 572351 215078 573151
rect 219162 572351 219218 573151
rect 223394 572351 223450 573151
rect 227534 572351 227590 573151
rect 231766 572351 231822 573151
rect 235906 572351 235962 573151
rect 240138 572351 240194 573151
rect 244278 572351 244334 573151
rect 248418 572351 248474 573151
rect 252650 572351 252706 573151
rect 256790 572351 256846 573151
rect 261022 572351 261078 573151
rect 265162 572351 265218 573151
rect 269302 572351 269358 573151
rect 273534 572351 273590 573151
rect 277674 572351 277730 573151
rect 281906 572351 281962 573151
rect 286046 572351 286102 573151
rect 290186 572351 290242 573151
rect 294418 572351 294474 573151
rect 298558 572351 298614 573151
rect 302790 572351 302846 573151
rect 306930 572351 306986 573151
rect 311070 572351 311126 573151
rect 315302 572351 315358 573151
rect 319442 572351 319498 573151
rect 323674 572351 323730 573151
rect 327814 572351 327870 573151
rect 331954 572351 332010 573151
rect 336186 572351 336242 573151
rect 340326 572351 340382 573151
rect 344558 572351 344614 573151
rect 348698 572351 348754 573151
rect 352838 572351 352894 573151
rect 357070 572351 357126 573151
rect 361210 572351 361266 573151
rect 365442 572351 365498 573151
rect 369582 572351 369638 573151
rect 373722 572351 373778 573151
rect 377954 572351 378010 573151
rect 382094 572351 382150 573151
rect 386326 572351 386382 573151
rect 390466 572351 390522 573151
rect 394606 572351 394662 573151
rect 398838 572351 398894 573151
rect 402978 572351 403034 573151
rect 407210 572351 407266 573151
rect 411350 572351 411406 573151
rect 415490 572351 415546 573151
rect 419722 572351 419778 573151
rect 423862 572351 423918 573151
rect 428094 572351 428150 573151
rect 432234 572351 432290 573151
rect 436374 572351 436430 573151
rect 440606 572351 440662 573151
rect 444746 572351 444802 573151
rect 448978 572351 449034 573151
rect 453118 572351 453174 573151
rect 457258 572351 457314 573151
rect 461490 572351 461546 573151
rect 465630 572351 465686 573151
rect 469862 572351 469918 573151
rect 474002 572351 474058 573151
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3330 0 3386 800
rect 4250 0 4306 800
rect 5262 0 5318 800
rect 6182 0 6238 800
rect 7194 0 7250 800
rect 8114 0 8170 800
rect 9126 0 9182 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12990 0 13046 800
rect 13910 0 13966 800
rect 14922 0 14978 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17774 0 17830 800
rect 18786 0 18842 800
rect 19706 0 19762 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22650 0 22706 800
rect 23570 0 23626 800
rect 24582 0 24638 800
rect 25502 0 25558 800
rect 26514 0 26570 800
rect 27434 0 27490 800
rect 28446 0 28502 800
rect 29366 0 29422 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 32310 0 32366 800
rect 33230 0 33286 800
rect 34242 0 34298 800
rect 35162 0 35218 800
rect 36174 0 36230 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39026 0 39082 800
rect 40038 0 40094 800
rect 40958 0 41014 800
rect 41970 0 42026 800
rect 42890 0 42946 800
rect 43902 0 43958 800
rect 44822 0 44878 800
rect 45834 0 45890 800
rect 46754 0 46810 800
rect 47766 0 47822 800
rect 48686 0 48742 800
rect 49698 0 49754 800
rect 50618 0 50674 800
rect 51630 0 51686 800
rect 52550 0 52606 800
rect 53562 0 53618 800
rect 54482 0 54538 800
rect 55494 0 55550 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60278 0 60334 800
rect 61290 0 61346 800
rect 62210 0 62266 800
rect 63222 0 63278 800
rect 64142 0 64198 800
rect 65154 0 65210 800
rect 66074 0 66130 800
rect 67086 0 67142 800
rect 68006 0 68062 800
rect 69018 0 69074 800
rect 69938 0 69994 800
rect 70950 0 71006 800
rect 71870 0 71926 800
rect 72882 0 72938 800
rect 73802 0 73858 800
rect 74814 0 74870 800
rect 75734 0 75790 800
rect 76746 0 76802 800
rect 77666 0 77722 800
rect 78678 0 78734 800
rect 79598 0 79654 800
rect 80610 0 80666 800
rect 81530 0 81586 800
rect 82542 0 82598 800
rect 83462 0 83518 800
rect 84474 0 84530 800
rect 85394 0 85450 800
rect 86406 0 86462 800
rect 87326 0 87382 800
rect 88338 0 88394 800
rect 89258 0 89314 800
rect 90270 0 90326 800
rect 91190 0 91246 800
rect 92202 0 92258 800
rect 93122 0 93178 800
rect 94134 0 94190 800
rect 95054 0 95110 800
rect 96066 0 96122 800
rect 96986 0 97042 800
rect 97998 0 98054 800
rect 98918 0 98974 800
rect 99930 0 99986 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102782 0 102838 800
rect 103794 0 103850 800
rect 104714 0 104770 800
rect 105726 0 105782 800
rect 106646 0 106702 800
rect 107658 0 107714 800
rect 108578 0 108634 800
rect 109590 0 109646 800
rect 110510 0 110566 800
rect 111522 0 111578 800
rect 112442 0 112498 800
rect 113454 0 113510 800
rect 114374 0 114430 800
rect 115386 0 115442 800
rect 116306 0 116362 800
rect 117318 0 117374 800
rect 118238 0 118294 800
rect 119250 0 119306 800
rect 120170 0 120226 800
rect 121182 0 121238 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124034 0 124090 800
rect 125046 0 125102 800
rect 125966 0 126022 800
rect 126978 0 127034 800
rect 127898 0 127954 800
rect 128910 0 128966 800
rect 129830 0 129886 800
rect 130842 0 130898 800
rect 131762 0 131818 800
rect 132774 0 132830 800
rect 133694 0 133750 800
rect 134706 0 134762 800
rect 135626 0 135682 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139490 0 139546 800
rect 140502 0 140558 800
rect 141422 0 141478 800
rect 142434 0 142490 800
rect 143354 0 143410 800
rect 144366 0 144422 800
rect 145286 0 145342 800
rect 146298 0 146354 800
rect 147218 0 147274 800
rect 148230 0 148286 800
rect 149150 0 149206 800
rect 150162 0 150218 800
rect 151082 0 151138 800
rect 152094 0 152150 800
rect 153014 0 153070 800
rect 154026 0 154082 800
rect 154946 0 155002 800
rect 155958 0 156014 800
rect 156878 0 156934 800
rect 157890 0 157946 800
rect 158810 0 158866 800
rect 159822 0 159878 800
rect 160742 0 160798 800
rect 161754 0 161810 800
rect 162674 0 162730 800
rect 163686 0 163742 800
rect 164606 0 164662 800
rect 165618 0 165674 800
rect 166538 0 166594 800
rect 167550 0 167606 800
rect 168470 0 168526 800
rect 169482 0 169538 800
rect 170402 0 170458 800
rect 171414 0 171470 800
rect 172334 0 172390 800
rect 173346 0 173402 800
rect 174266 0 174322 800
rect 175278 0 175334 800
rect 176198 0 176254 800
rect 177210 0 177266 800
rect 178130 0 178186 800
rect 179142 0 179198 800
rect 180062 0 180118 800
rect 181074 0 181130 800
rect 181994 0 182050 800
rect 183006 0 183062 800
rect 183926 0 183982 800
rect 184938 0 184994 800
rect 185858 0 185914 800
rect 186870 0 186926 800
rect 187790 0 187846 800
rect 188802 0 188858 800
rect 189722 0 189778 800
rect 190734 0 190790 800
rect 191654 0 191710 800
rect 192666 0 192722 800
rect 193586 0 193642 800
rect 194598 0 194654 800
rect 195518 0 195574 800
rect 196530 0 196586 800
rect 197450 0 197506 800
rect 198462 0 198518 800
rect 199382 0 199438 800
rect 200394 0 200450 800
rect 201314 0 201370 800
rect 202326 0 202382 800
rect 203246 0 203302 800
rect 204258 0 204314 800
rect 205178 0 205234 800
rect 206190 0 206246 800
rect 207110 0 207166 800
rect 208122 0 208178 800
rect 209042 0 209098 800
rect 210054 0 210110 800
rect 210974 0 211030 800
rect 211986 0 212042 800
rect 212906 0 212962 800
rect 213918 0 213974 800
rect 214838 0 214894 800
rect 215850 0 215906 800
rect 216770 0 216826 800
rect 217782 0 217838 800
rect 218702 0 218758 800
rect 219714 0 219770 800
rect 220634 0 220690 800
rect 221646 0 221702 800
rect 222566 0 222622 800
rect 223578 0 223634 800
rect 224498 0 224554 800
rect 225510 0 225566 800
rect 226430 0 226486 800
rect 227442 0 227498 800
rect 228362 0 228418 800
rect 229374 0 229430 800
rect 230294 0 230350 800
rect 231306 0 231362 800
rect 232226 0 232282 800
rect 233238 0 233294 800
rect 234158 0 234214 800
rect 235170 0 235226 800
rect 236090 0 236146 800
rect 237102 0 237158 800
rect 238022 0 238078 800
rect 239034 0 239090 800
rect 239954 0 240010 800
rect 240966 0 241022 800
rect 241886 0 241942 800
rect 242898 0 242954 800
rect 243818 0 243874 800
rect 244830 0 244886 800
rect 245750 0 245806 800
rect 246762 0 246818 800
rect 247682 0 247738 800
rect 248694 0 248750 800
rect 249614 0 249670 800
rect 250626 0 250682 800
rect 251546 0 251602 800
rect 252558 0 252614 800
rect 253478 0 253534 800
rect 254490 0 254546 800
rect 255410 0 255466 800
rect 256422 0 256478 800
rect 257342 0 257398 800
rect 258354 0 258410 800
rect 259274 0 259330 800
rect 260286 0 260342 800
rect 261206 0 261262 800
rect 262218 0 262274 800
rect 263138 0 263194 800
rect 264150 0 264206 800
rect 265070 0 265126 800
rect 266082 0 266138 800
rect 267002 0 267058 800
rect 268014 0 268070 800
rect 268934 0 268990 800
rect 269946 0 270002 800
rect 270866 0 270922 800
rect 271878 0 271934 800
rect 272798 0 272854 800
rect 273810 0 273866 800
rect 274730 0 274786 800
rect 275742 0 275798 800
rect 276662 0 276718 800
rect 277674 0 277730 800
rect 278594 0 278650 800
rect 279606 0 279662 800
rect 280526 0 280582 800
rect 281538 0 281594 800
rect 282458 0 282514 800
rect 283470 0 283526 800
rect 284390 0 284446 800
rect 285402 0 285458 800
rect 286322 0 286378 800
rect 287334 0 287390 800
rect 288254 0 288310 800
rect 289266 0 289322 800
rect 290186 0 290242 800
rect 291198 0 291254 800
rect 292118 0 292174 800
rect 293130 0 293186 800
rect 294050 0 294106 800
rect 295062 0 295118 800
rect 295982 0 296038 800
rect 296994 0 297050 800
rect 297914 0 297970 800
rect 298926 0 298982 800
rect 299846 0 299902 800
rect 300858 0 300914 800
rect 301778 0 301834 800
rect 302790 0 302846 800
rect 303710 0 303766 800
rect 304722 0 304778 800
rect 305642 0 305698 800
rect 306654 0 306710 800
rect 307574 0 307630 800
rect 308586 0 308642 800
rect 309506 0 309562 800
rect 310518 0 310574 800
rect 311438 0 311494 800
rect 312450 0 312506 800
rect 313370 0 313426 800
rect 314382 0 314438 800
rect 315302 0 315358 800
rect 316314 0 316370 800
rect 317234 0 317290 800
rect 318246 0 318302 800
rect 319166 0 319222 800
rect 320178 0 320234 800
rect 321098 0 321154 800
rect 322110 0 322166 800
rect 323030 0 323086 800
rect 324042 0 324098 800
rect 324962 0 325018 800
rect 325974 0 326030 800
rect 326894 0 326950 800
rect 327906 0 327962 800
rect 328826 0 328882 800
rect 329838 0 329894 800
rect 330758 0 330814 800
rect 331770 0 331826 800
rect 332690 0 332746 800
rect 333702 0 333758 800
rect 334622 0 334678 800
rect 335634 0 335690 800
rect 336554 0 336610 800
rect 337566 0 337622 800
rect 338486 0 338542 800
rect 339498 0 339554 800
rect 340418 0 340474 800
rect 341430 0 341486 800
rect 342350 0 342406 800
rect 343362 0 343418 800
rect 344282 0 344338 800
rect 345294 0 345350 800
rect 346214 0 346270 800
rect 347226 0 347282 800
rect 348146 0 348202 800
rect 349158 0 349214 800
rect 350078 0 350134 800
rect 351090 0 351146 800
rect 352010 0 352066 800
rect 353022 0 353078 800
rect 353942 0 353998 800
rect 354954 0 355010 800
rect 355874 0 355930 800
rect 356886 0 356942 800
rect 357806 0 357862 800
rect 358818 0 358874 800
rect 359738 0 359794 800
rect 360750 0 360806 800
rect 361670 0 361726 800
rect 362682 0 362738 800
rect 363602 0 363658 800
rect 364614 0 364670 800
rect 365534 0 365590 800
rect 366546 0 366602 800
rect 367466 0 367522 800
rect 368478 0 368534 800
rect 369398 0 369454 800
rect 370410 0 370466 800
rect 371330 0 371386 800
rect 372342 0 372398 800
rect 373262 0 373318 800
rect 374274 0 374330 800
rect 375194 0 375250 800
rect 376206 0 376262 800
rect 377126 0 377182 800
rect 378138 0 378194 800
rect 379058 0 379114 800
rect 380070 0 380126 800
rect 380990 0 381046 800
rect 382002 0 382058 800
rect 382922 0 382978 800
rect 383934 0 383990 800
rect 384854 0 384910 800
rect 385866 0 385922 800
rect 386786 0 386842 800
rect 387798 0 387854 800
rect 388718 0 388774 800
rect 389730 0 389786 800
rect 390650 0 390706 800
rect 391662 0 391718 800
rect 392582 0 392638 800
rect 393594 0 393650 800
rect 394514 0 394570 800
rect 395526 0 395582 800
rect 396446 0 396502 800
rect 397458 0 397514 800
rect 398378 0 398434 800
rect 399390 0 399446 800
rect 400310 0 400366 800
rect 401322 0 401378 800
rect 402242 0 402298 800
rect 403254 0 403310 800
rect 404174 0 404230 800
rect 405186 0 405242 800
rect 406106 0 406162 800
rect 407118 0 407174 800
rect 408038 0 408094 800
rect 409050 0 409106 800
rect 409970 0 410026 800
rect 410982 0 411038 800
rect 411902 0 411958 800
rect 412914 0 412970 800
rect 413834 0 413890 800
rect 414846 0 414902 800
rect 415766 0 415822 800
rect 416778 0 416834 800
rect 417698 0 417754 800
rect 418710 0 418766 800
rect 419630 0 419686 800
rect 420642 0 420698 800
rect 421562 0 421618 800
rect 422574 0 422630 800
rect 423494 0 423550 800
rect 424506 0 424562 800
rect 425426 0 425482 800
rect 426438 0 426494 800
rect 427358 0 427414 800
rect 428370 0 428426 800
rect 429290 0 429346 800
rect 430302 0 430358 800
rect 431222 0 431278 800
rect 432234 0 432290 800
rect 433154 0 433210 800
rect 434166 0 434222 800
rect 435086 0 435142 800
rect 436098 0 436154 800
rect 437018 0 437074 800
rect 438030 0 438086 800
rect 438950 0 439006 800
rect 439962 0 440018 800
rect 440882 0 440938 800
rect 441894 0 441950 800
rect 442814 0 442870 800
rect 443826 0 443882 800
rect 444746 0 444802 800
rect 445758 0 445814 800
rect 446678 0 446734 800
rect 447690 0 447746 800
rect 448610 0 448666 800
rect 449622 0 449678 800
rect 450542 0 450598 800
rect 451554 0 451610 800
rect 452474 0 452530 800
rect 453486 0 453542 800
rect 454406 0 454462 800
rect 455418 0 455474 800
rect 456338 0 456394 800
rect 457350 0 457406 800
rect 458270 0 458326 800
rect 459282 0 459338 800
rect 460202 0 460258 800
rect 461214 0 461270 800
rect 462134 0 462190 800
rect 463146 0 463202 800
rect 464066 0 464122 800
rect 465078 0 465134 800
rect 465998 0 466054 800
rect 467010 0 467066 800
rect 467930 0 467986 800
rect 468942 0 468998 800
rect 469862 0 469918 800
rect 470874 0 470930 800
rect 471794 0 471850 800
rect 472806 0 472862 800
rect 473726 0 473782 800
rect 474738 0 474794 800
rect 475658 0 475714 800
<< obsm2 >>
rect 480 572295 1986 572351
rect 2154 572295 6126 572351
rect 6294 572295 10266 572351
rect 10434 572295 14498 572351
rect 14666 572295 18638 572351
rect 18806 572295 22870 572351
rect 23038 572295 27010 572351
rect 27178 572295 31150 572351
rect 31318 572295 35382 572351
rect 35550 572295 39522 572351
rect 39690 572295 43754 572351
rect 43922 572295 47894 572351
rect 48062 572295 52034 572351
rect 52202 572295 56266 572351
rect 56434 572295 60406 572351
rect 60574 572295 64638 572351
rect 64806 572295 68778 572351
rect 68946 572295 72918 572351
rect 73086 572295 77150 572351
rect 77318 572295 81290 572351
rect 81458 572295 85522 572351
rect 85690 572295 89662 572351
rect 89830 572295 93802 572351
rect 93970 572295 98034 572351
rect 98202 572295 102174 572351
rect 102342 572295 106406 572351
rect 106574 572295 110546 572351
rect 110714 572295 114686 572351
rect 114854 572295 118918 572351
rect 119086 572295 123058 572351
rect 123226 572295 127290 572351
rect 127458 572295 131430 572351
rect 131598 572295 135570 572351
rect 135738 572295 139802 572351
rect 139970 572295 143942 572351
rect 144110 572295 148174 572351
rect 148342 572295 152314 572351
rect 152482 572295 156454 572351
rect 156622 572295 160686 572351
rect 160854 572295 164826 572351
rect 164994 572295 169058 572351
rect 169226 572295 173198 572351
rect 173366 572295 177338 572351
rect 177506 572295 181570 572351
rect 181738 572295 185710 572351
rect 185878 572295 189942 572351
rect 190110 572295 194082 572351
rect 194250 572295 198222 572351
rect 198390 572295 202454 572351
rect 202622 572295 206594 572351
rect 206762 572295 210826 572351
rect 210994 572295 214966 572351
rect 215134 572295 219106 572351
rect 219274 572295 223338 572351
rect 223506 572295 227478 572351
rect 227646 572295 231710 572351
rect 231878 572295 235850 572351
rect 236018 572295 240082 572351
rect 240250 572295 244222 572351
rect 244390 572295 248362 572351
rect 248530 572295 252594 572351
rect 252762 572295 256734 572351
rect 256902 572295 260966 572351
rect 261134 572295 265106 572351
rect 265274 572295 269246 572351
rect 269414 572295 273478 572351
rect 273646 572295 277618 572351
rect 277786 572295 281850 572351
rect 282018 572295 285990 572351
rect 286158 572295 290130 572351
rect 290298 572295 294362 572351
rect 294530 572295 298502 572351
rect 298670 572295 302734 572351
rect 302902 572295 306874 572351
rect 307042 572295 311014 572351
rect 311182 572295 315246 572351
rect 315414 572295 319386 572351
rect 319554 572295 323618 572351
rect 323786 572295 327758 572351
rect 327926 572295 331898 572351
rect 332066 572295 336130 572351
rect 336298 572295 340270 572351
rect 340438 572295 344502 572351
rect 344670 572295 348642 572351
rect 348810 572295 352782 572351
rect 352950 572295 357014 572351
rect 357182 572295 361154 572351
rect 361322 572295 365386 572351
rect 365554 572295 369526 572351
rect 369694 572295 373666 572351
rect 373834 572295 377898 572351
rect 378066 572295 382038 572351
rect 382206 572295 386270 572351
rect 386438 572295 390410 572351
rect 390578 572295 394550 572351
rect 394718 572295 398782 572351
rect 398950 572295 402922 572351
rect 403090 572295 407154 572351
rect 407322 572295 411294 572351
rect 411462 572295 415434 572351
rect 415602 572295 419666 572351
rect 419834 572295 423806 572351
rect 423974 572295 428038 572351
rect 428206 572295 432178 572351
rect 432346 572295 436318 572351
rect 436486 572295 440550 572351
rect 440718 572295 444690 572351
rect 444858 572295 448922 572351
rect 449090 572295 453062 572351
rect 453230 572295 457202 572351
rect 457370 572295 461434 572351
rect 461602 572295 465574 572351
rect 465742 572295 469806 572351
rect 469974 572295 473946 572351
rect 474114 572295 475712 572351
rect 480 856 475712 572295
rect 590 2 1342 856
rect 1510 2 2262 856
rect 2430 2 3274 856
rect 3442 2 4194 856
rect 4362 2 5206 856
rect 5374 2 6126 856
rect 6294 2 7138 856
rect 7306 2 8058 856
rect 8226 2 9070 856
rect 9238 2 9990 856
rect 10158 2 11002 856
rect 11170 2 11922 856
rect 12090 2 12934 856
rect 13102 2 13854 856
rect 14022 2 14866 856
rect 15034 2 15786 856
rect 15954 2 16798 856
rect 16966 2 17718 856
rect 17886 2 18730 856
rect 18898 2 19650 856
rect 19818 2 20662 856
rect 20830 2 21582 856
rect 21750 2 22594 856
rect 22762 2 23514 856
rect 23682 2 24526 856
rect 24694 2 25446 856
rect 25614 2 26458 856
rect 26626 2 27378 856
rect 27546 2 28390 856
rect 28558 2 29310 856
rect 29478 2 30322 856
rect 30490 2 31242 856
rect 31410 2 32254 856
rect 32422 2 33174 856
rect 33342 2 34186 856
rect 34354 2 35106 856
rect 35274 2 36118 856
rect 36286 2 37038 856
rect 37206 2 38050 856
rect 38218 2 38970 856
rect 39138 2 39982 856
rect 40150 2 40902 856
rect 41070 2 41914 856
rect 42082 2 42834 856
rect 43002 2 43846 856
rect 44014 2 44766 856
rect 44934 2 45778 856
rect 45946 2 46698 856
rect 46866 2 47710 856
rect 47878 2 48630 856
rect 48798 2 49642 856
rect 49810 2 50562 856
rect 50730 2 51574 856
rect 51742 2 52494 856
rect 52662 2 53506 856
rect 53674 2 54426 856
rect 54594 2 55438 856
rect 55606 2 56358 856
rect 56526 2 57370 856
rect 57538 2 58290 856
rect 58458 2 59302 856
rect 59470 2 60222 856
rect 60390 2 61234 856
rect 61402 2 62154 856
rect 62322 2 63166 856
rect 63334 2 64086 856
rect 64254 2 65098 856
rect 65266 2 66018 856
rect 66186 2 67030 856
rect 67198 2 67950 856
rect 68118 2 68962 856
rect 69130 2 69882 856
rect 70050 2 70894 856
rect 71062 2 71814 856
rect 71982 2 72826 856
rect 72994 2 73746 856
rect 73914 2 74758 856
rect 74926 2 75678 856
rect 75846 2 76690 856
rect 76858 2 77610 856
rect 77778 2 78622 856
rect 78790 2 79542 856
rect 79710 2 80554 856
rect 80722 2 81474 856
rect 81642 2 82486 856
rect 82654 2 83406 856
rect 83574 2 84418 856
rect 84586 2 85338 856
rect 85506 2 86350 856
rect 86518 2 87270 856
rect 87438 2 88282 856
rect 88450 2 89202 856
rect 89370 2 90214 856
rect 90382 2 91134 856
rect 91302 2 92146 856
rect 92314 2 93066 856
rect 93234 2 94078 856
rect 94246 2 94998 856
rect 95166 2 96010 856
rect 96178 2 96930 856
rect 97098 2 97942 856
rect 98110 2 98862 856
rect 99030 2 99874 856
rect 100042 2 100794 856
rect 100962 2 101806 856
rect 101974 2 102726 856
rect 102894 2 103738 856
rect 103906 2 104658 856
rect 104826 2 105670 856
rect 105838 2 106590 856
rect 106758 2 107602 856
rect 107770 2 108522 856
rect 108690 2 109534 856
rect 109702 2 110454 856
rect 110622 2 111466 856
rect 111634 2 112386 856
rect 112554 2 113398 856
rect 113566 2 114318 856
rect 114486 2 115330 856
rect 115498 2 116250 856
rect 116418 2 117262 856
rect 117430 2 118182 856
rect 118350 2 119194 856
rect 119362 2 120114 856
rect 120282 2 121126 856
rect 121294 2 122046 856
rect 122214 2 123058 856
rect 123226 2 123978 856
rect 124146 2 124990 856
rect 125158 2 125910 856
rect 126078 2 126922 856
rect 127090 2 127842 856
rect 128010 2 128854 856
rect 129022 2 129774 856
rect 129942 2 130786 856
rect 130954 2 131706 856
rect 131874 2 132718 856
rect 132886 2 133638 856
rect 133806 2 134650 856
rect 134818 2 135570 856
rect 135738 2 136582 856
rect 136750 2 137502 856
rect 137670 2 138514 856
rect 138682 2 139434 856
rect 139602 2 140446 856
rect 140614 2 141366 856
rect 141534 2 142378 856
rect 142546 2 143298 856
rect 143466 2 144310 856
rect 144478 2 145230 856
rect 145398 2 146242 856
rect 146410 2 147162 856
rect 147330 2 148174 856
rect 148342 2 149094 856
rect 149262 2 150106 856
rect 150274 2 151026 856
rect 151194 2 152038 856
rect 152206 2 152958 856
rect 153126 2 153970 856
rect 154138 2 154890 856
rect 155058 2 155902 856
rect 156070 2 156822 856
rect 156990 2 157834 856
rect 158002 2 158754 856
rect 158922 2 159766 856
rect 159934 2 160686 856
rect 160854 2 161698 856
rect 161866 2 162618 856
rect 162786 2 163630 856
rect 163798 2 164550 856
rect 164718 2 165562 856
rect 165730 2 166482 856
rect 166650 2 167494 856
rect 167662 2 168414 856
rect 168582 2 169426 856
rect 169594 2 170346 856
rect 170514 2 171358 856
rect 171526 2 172278 856
rect 172446 2 173290 856
rect 173458 2 174210 856
rect 174378 2 175222 856
rect 175390 2 176142 856
rect 176310 2 177154 856
rect 177322 2 178074 856
rect 178242 2 179086 856
rect 179254 2 180006 856
rect 180174 2 181018 856
rect 181186 2 181938 856
rect 182106 2 182950 856
rect 183118 2 183870 856
rect 184038 2 184882 856
rect 185050 2 185802 856
rect 185970 2 186814 856
rect 186982 2 187734 856
rect 187902 2 188746 856
rect 188914 2 189666 856
rect 189834 2 190678 856
rect 190846 2 191598 856
rect 191766 2 192610 856
rect 192778 2 193530 856
rect 193698 2 194542 856
rect 194710 2 195462 856
rect 195630 2 196474 856
rect 196642 2 197394 856
rect 197562 2 198406 856
rect 198574 2 199326 856
rect 199494 2 200338 856
rect 200506 2 201258 856
rect 201426 2 202270 856
rect 202438 2 203190 856
rect 203358 2 204202 856
rect 204370 2 205122 856
rect 205290 2 206134 856
rect 206302 2 207054 856
rect 207222 2 208066 856
rect 208234 2 208986 856
rect 209154 2 209998 856
rect 210166 2 210918 856
rect 211086 2 211930 856
rect 212098 2 212850 856
rect 213018 2 213862 856
rect 214030 2 214782 856
rect 214950 2 215794 856
rect 215962 2 216714 856
rect 216882 2 217726 856
rect 217894 2 218646 856
rect 218814 2 219658 856
rect 219826 2 220578 856
rect 220746 2 221590 856
rect 221758 2 222510 856
rect 222678 2 223522 856
rect 223690 2 224442 856
rect 224610 2 225454 856
rect 225622 2 226374 856
rect 226542 2 227386 856
rect 227554 2 228306 856
rect 228474 2 229318 856
rect 229486 2 230238 856
rect 230406 2 231250 856
rect 231418 2 232170 856
rect 232338 2 233182 856
rect 233350 2 234102 856
rect 234270 2 235114 856
rect 235282 2 236034 856
rect 236202 2 237046 856
rect 237214 2 237966 856
rect 238134 2 238978 856
rect 239146 2 239898 856
rect 240066 2 240910 856
rect 241078 2 241830 856
rect 241998 2 242842 856
rect 243010 2 243762 856
rect 243930 2 244774 856
rect 244942 2 245694 856
rect 245862 2 246706 856
rect 246874 2 247626 856
rect 247794 2 248638 856
rect 248806 2 249558 856
rect 249726 2 250570 856
rect 250738 2 251490 856
rect 251658 2 252502 856
rect 252670 2 253422 856
rect 253590 2 254434 856
rect 254602 2 255354 856
rect 255522 2 256366 856
rect 256534 2 257286 856
rect 257454 2 258298 856
rect 258466 2 259218 856
rect 259386 2 260230 856
rect 260398 2 261150 856
rect 261318 2 262162 856
rect 262330 2 263082 856
rect 263250 2 264094 856
rect 264262 2 265014 856
rect 265182 2 266026 856
rect 266194 2 266946 856
rect 267114 2 267958 856
rect 268126 2 268878 856
rect 269046 2 269890 856
rect 270058 2 270810 856
rect 270978 2 271822 856
rect 271990 2 272742 856
rect 272910 2 273754 856
rect 273922 2 274674 856
rect 274842 2 275686 856
rect 275854 2 276606 856
rect 276774 2 277618 856
rect 277786 2 278538 856
rect 278706 2 279550 856
rect 279718 2 280470 856
rect 280638 2 281482 856
rect 281650 2 282402 856
rect 282570 2 283414 856
rect 283582 2 284334 856
rect 284502 2 285346 856
rect 285514 2 286266 856
rect 286434 2 287278 856
rect 287446 2 288198 856
rect 288366 2 289210 856
rect 289378 2 290130 856
rect 290298 2 291142 856
rect 291310 2 292062 856
rect 292230 2 293074 856
rect 293242 2 293994 856
rect 294162 2 295006 856
rect 295174 2 295926 856
rect 296094 2 296938 856
rect 297106 2 297858 856
rect 298026 2 298870 856
rect 299038 2 299790 856
rect 299958 2 300802 856
rect 300970 2 301722 856
rect 301890 2 302734 856
rect 302902 2 303654 856
rect 303822 2 304666 856
rect 304834 2 305586 856
rect 305754 2 306598 856
rect 306766 2 307518 856
rect 307686 2 308530 856
rect 308698 2 309450 856
rect 309618 2 310462 856
rect 310630 2 311382 856
rect 311550 2 312394 856
rect 312562 2 313314 856
rect 313482 2 314326 856
rect 314494 2 315246 856
rect 315414 2 316258 856
rect 316426 2 317178 856
rect 317346 2 318190 856
rect 318358 2 319110 856
rect 319278 2 320122 856
rect 320290 2 321042 856
rect 321210 2 322054 856
rect 322222 2 322974 856
rect 323142 2 323986 856
rect 324154 2 324906 856
rect 325074 2 325918 856
rect 326086 2 326838 856
rect 327006 2 327850 856
rect 328018 2 328770 856
rect 328938 2 329782 856
rect 329950 2 330702 856
rect 330870 2 331714 856
rect 331882 2 332634 856
rect 332802 2 333646 856
rect 333814 2 334566 856
rect 334734 2 335578 856
rect 335746 2 336498 856
rect 336666 2 337510 856
rect 337678 2 338430 856
rect 338598 2 339442 856
rect 339610 2 340362 856
rect 340530 2 341374 856
rect 341542 2 342294 856
rect 342462 2 343306 856
rect 343474 2 344226 856
rect 344394 2 345238 856
rect 345406 2 346158 856
rect 346326 2 347170 856
rect 347338 2 348090 856
rect 348258 2 349102 856
rect 349270 2 350022 856
rect 350190 2 351034 856
rect 351202 2 351954 856
rect 352122 2 352966 856
rect 353134 2 353886 856
rect 354054 2 354898 856
rect 355066 2 355818 856
rect 355986 2 356830 856
rect 356998 2 357750 856
rect 357918 2 358762 856
rect 358930 2 359682 856
rect 359850 2 360694 856
rect 360862 2 361614 856
rect 361782 2 362626 856
rect 362794 2 363546 856
rect 363714 2 364558 856
rect 364726 2 365478 856
rect 365646 2 366490 856
rect 366658 2 367410 856
rect 367578 2 368422 856
rect 368590 2 369342 856
rect 369510 2 370354 856
rect 370522 2 371274 856
rect 371442 2 372286 856
rect 372454 2 373206 856
rect 373374 2 374218 856
rect 374386 2 375138 856
rect 375306 2 376150 856
rect 376318 2 377070 856
rect 377238 2 378082 856
rect 378250 2 379002 856
rect 379170 2 380014 856
rect 380182 2 380934 856
rect 381102 2 381946 856
rect 382114 2 382866 856
rect 383034 2 383878 856
rect 384046 2 384798 856
rect 384966 2 385810 856
rect 385978 2 386730 856
rect 386898 2 387742 856
rect 387910 2 388662 856
rect 388830 2 389674 856
rect 389842 2 390594 856
rect 390762 2 391606 856
rect 391774 2 392526 856
rect 392694 2 393538 856
rect 393706 2 394458 856
rect 394626 2 395470 856
rect 395638 2 396390 856
rect 396558 2 397402 856
rect 397570 2 398322 856
rect 398490 2 399334 856
rect 399502 2 400254 856
rect 400422 2 401266 856
rect 401434 2 402186 856
rect 402354 2 403198 856
rect 403366 2 404118 856
rect 404286 2 405130 856
rect 405298 2 406050 856
rect 406218 2 407062 856
rect 407230 2 407982 856
rect 408150 2 408994 856
rect 409162 2 409914 856
rect 410082 2 410926 856
rect 411094 2 411846 856
rect 412014 2 412858 856
rect 413026 2 413778 856
rect 413946 2 414790 856
rect 414958 2 415710 856
rect 415878 2 416722 856
rect 416890 2 417642 856
rect 417810 2 418654 856
rect 418822 2 419574 856
rect 419742 2 420586 856
rect 420754 2 421506 856
rect 421674 2 422518 856
rect 422686 2 423438 856
rect 423606 2 424450 856
rect 424618 2 425370 856
rect 425538 2 426382 856
rect 426550 2 427302 856
rect 427470 2 428314 856
rect 428482 2 429234 856
rect 429402 2 430246 856
rect 430414 2 431166 856
rect 431334 2 432178 856
rect 432346 2 433098 856
rect 433266 2 434110 856
rect 434278 2 435030 856
rect 435198 2 436042 856
rect 436210 2 436962 856
rect 437130 2 437974 856
rect 438142 2 438894 856
rect 439062 2 439906 856
rect 440074 2 440826 856
rect 440994 2 441838 856
rect 442006 2 442758 856
rect 442926 2 443770 856
rect 443938 2 444690 856
rect 444858 2 445702 856
rect 445870 2 446622 856
rect 446790 2 447634 856
rect 447802 2 448554 856
rect 448722 2 449566 856
rect 449734 2 450486 856
rect 450654 2 451498 856
rect 451666 2 452418 856
rect 452586 2 453430 856
rect 453598 2 454350 856
rect 454518 2 455362 856
rect 455530 2 456282 856
rect 456450 2 457294 856
rect 457462 2 458214 856
rect 458382 2 459226 856
rect 459394 2 460146 856
rect 460314 2 461158 856
rect 461326 2 462078 856
rect 462246 2 463090 856
rect 463258 2 464010 856
rect 464178 2 465022 856
rect 465190 2 465942 856
rect 466110 2 466954 856
rect 467122 2 467874 856
rect 468042 2 468886 856
rect 469054 2 469806 856
rect 469974 2 470818 856
rect 470986 2 471738 856
rect 471906 2 472750 856
rect 472918 2 473670 856
rect 473838 2 474682 856
rect 474850 2 475602 856
<< obsm3 >>
rect 2957 715 473235 570689
<< metal4 >>
rect 4208 2128 4528 570704
rect 19568 2128 19888 570704
rect 34928 2128 35248 570704
rect 50288 2128 50608 570704
rect 65648 2128 65968 570704
rect 81008 2128 81328 570704
rect 96368 2128 96688 570704
rect 111728 2128 112048 570704
rect 127088 2128 127408 570704
rect 142448 2128 142768 570704
rect 157808 2128 158128 570704
rect 173168 2128 173488 570704
rect 188528 2128 188848 570704
rect 203888 2128 204208 570704
rect 219248 2128 219568 570704
rect 234608 2128 234928 570704
rect 249968 2128 250288 570704
rect 265328 2128 265648 570704
rect 280688 2128 281008 570704
rect 296048 2128 296368 570704
rect 311408 2128 311728 570704
rect 326768 2128 327088 570704
rect 342128 2128 342448 570704
rect 357488 2128 357808 570704
rect 372848 2128 373168 570704
rect 388208 2128 388528 570704
rect 403568 2128 403888 570704
rect 418928 2128 419248 570704
rect 434288 2128 434608 570704
rect 449648 2128 449968 570704
rect 465008 2128 465328 570704
<< obsm4 >>
rect 18827 2755 19488 550357
rect 19968 2755 34848 550357
rect 35328 2755 50208 550357
rect 50688 2755 65568 550357
rect 66048 2755 80928 550357
rect 81408 2755 96288 550357
rect 96768 2755 111648 550357
rect 112128 2755 127008 550357
rect 127488 2755 142368 550357
rect 142848 2755 157728 550357
rect 158208 2755 173088 550357
rect 173568 2755 188448 550357
rect 188928 2755 203808 550357
rect 204288 2755 219168 550357
rect 219648 2755 234528 550357
rect 235008 2755 249888 550357
rect 250368 2755 265248 550357
rect 265728 2755 280608 550357
rect 281088 2755 295968 550357
rect 296448 2755 311328 550357
rect 311808 2755 326688 550357
rect 327168 2755 342048 550357
rect 342528 2755 357408 550357
rect 357888 2755 372768 550357
rect 373248 2755 388128 550357
rect 388608 2755 403488 550357
rect 403968 2755 418848 550357
rect 419328 2755 434208 550357
rect 434688 2755 449568 550357
rect 450048 2755 464928 550357
rect 465408 2755 469141 550357
<< labels >>
rlabel metal2 s 2042 572351 2098 573151 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 127346 572351 127402 573151 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 139858 572351 139914 573151 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 152370 572351 152426 573151 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 164882 572351 164938 573151 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 177394 572351 177450 573151 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 189998 572351 190054 573151 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 202510 572351 202566 573151 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 215022 572351 215078 573151 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 227534 572351 227590 573151 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 240138 572351 240194 573151 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 14554 572351 14610 573151 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 252650 572351 252706 573151 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 265162 572351 265218 573151 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 277674 572351 277730 573151 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 290186 572351 290242 573151 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 302790 572351 302846 573151 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 315302 572351 315358 573151 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 327814 572351 327870 573151 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 340326 572351 340382 573151 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 352838 572351 352894 573151 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 365442 572351 365498 573151 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 27066 572351 27122 573151 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 377954 572351 378010 573151 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 390466 572351 390522 573151 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 402978 572351 403034 573151 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 415490 572351 415546 573151 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 428094 572351 428150 573151 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 440606 572351 440662 573151 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 453118 572351 453174 573151 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 465630 572351 465686 573151 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 39578 572351 39634 573151 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 52090 572351 52146 573151 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 64694 572351 64750 573151 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 77206 572351 77262 573151 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 89718 572351 89774 573151 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 102230 572351 102286 573151 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 114742 572351 114798 573151 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6182 572351 6238 573151 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 131486 572351 131542 573151 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 143998 572351 144054 573151 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 156510 572351 156566 573151 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 169114 572351 169170 573151 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 181626 572351 181682 573151 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 194138 572351 194194 573151 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 206650 572351 206706 573151 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 219162 572351 219218 573151 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 231766 572351 231822 573151 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 244278 572351 244334 573151 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 18694 572351 18750 573151 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 256790 572351 256846 573151 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 269302 572351 269358 573151 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 281906 572351 281962 573151 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 294418 572351 294474 573151 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 306930 572351 306986 573151 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 319442 572351 319498 573151 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 331954 572351 332010 573151 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 344558 572351 344614 573151 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 357070 572351 357126 573151 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 369582 572351 369638 573151 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 31206 572351 31262 573151 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 382094 572351 382150 573151 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 394606 572351 394662 573151 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 407210 572351 407266 573151 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 419722 572351 419778 573151 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 432234 572351 432290 573151 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 444746 572351 444802 573151 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 457258 572351 457314 573151 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 469862 572351 469918 573151 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 43810 572351 43866 573151 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 56322 572351 56378 573151 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 68834 572351 68890 573151 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 81346 572351 81402 573151 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 93858 572351 93914 573151 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 106462 572351 106518 573151 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 118974 572351 119030 573151 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 10322 572351 10378 573151 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 135626 572351 135682 573151 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 148230 572351 148286 573151 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 160742 572351 160798 573151 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 173254 572351 173310 573151 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 185766 572351 185822 573151 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 198278 572351 198334 573151 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 210882 572351 210938 573151 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 223394 572351 223450 573151 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 235906 572351 235962 573151 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 248418 572351 248474 573151 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 22926 572351 22982 573151 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 261022 572351 261078 573151 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 273534 572351 273590 573151 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 286046 572351 286102 573151 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 298558 572351 298614 573151 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 311070 572351 311126 573151 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 323674 572351 323730 573151 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 336186 572351 336242 573151 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 348698 572351 348754 573151 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 361210 572351 361266 573151 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 373722 572351 373778 573151 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 35438 572351 35494 573151 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 386326 572351 386382 573151 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 398838 572351 398894 573151 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 411350 572351 411406 573151 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 423862 572351 423918 573151 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 436374 572351 436430 573151 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 448978 572351 449034 573151 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 461490 572351 461546 573151 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 474002 572351 474058 573151 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 47950 572351 48006 573151 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 60462 572351 60518 573151 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 72974 572351 73030 573151 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 85578 572351 85634 573151 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 98090 572351 98146 573151 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 110602 572351 110658 573151 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 123114 572351 123170 573151 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 473726 0 473782 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 474738 0 474794 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 475658 0 475714 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 392582 0 392638 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 395526 0 395582 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 398378 0 398434 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 404174 0 404230 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 407118 0 407174 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 409970 0 410026 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 412914 0 412970 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 415766 0 415822 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 418710 0 418766 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 421562 0 421618 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 424506 0 424562 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 427358 0 427414 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 430302 0 430358 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 433154 0 433210 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 436098 0 436154 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 438950 0 439006 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 441894 0 441950 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 444746 0 444802 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 447690 0 447746 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 450542 0 450598 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 453486 0 453542 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 456338 0 456394 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 459282 0 459338 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 462134 0 462190 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 465078 0 465134 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 467930 0 467986 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 470874 0 470930 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 247682 0 247738 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 265070 0 265126 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 268014 0 268070 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 273810 0 273866 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 288254 0 288310 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 291198 0 291254 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 294050 0 294106 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 299846 0 299902 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 305642 0 305698 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 311438 0 311494 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 325974 0 326030 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 328826 0 328882 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 331770 0 331826 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 334622 0 334678 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 337566 0 337622 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 340418 0 340474 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 343362 0 343418 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 352010 0 352066 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 357806 0 357862 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 360750 0 360806 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 363602 0 363658 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 366546 0 366602 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 369398 0 369454 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 375194 0 375250 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 378138 0 378194 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 380990 0 381046 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 383934 0 383990 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 386786 0 386842 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 389730 0 389786 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 393594 0 393650 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 396446 0 396502 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 399390 0 399446 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 402242 0 402298 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 405186 0 405242 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 408038 0 408094 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 410982 0 411038 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 413834 0 413890 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 416778 0 416834 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 419630 0 419686 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 422574 0 422630 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 425426 0 425482 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 428370 0 428426 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 431222 0 431278 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 434166 0 434222 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 437018 0 437074 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 439962 0 440018 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 442814 0 442870 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 445758 0 445814 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 448610 0 448666 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 451554 0 451610 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 454406 0 454462 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 457350 0 457406 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 460202 0 460258 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 463146 0 463202 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 465998 0 466054 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 468942 0 468998 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 471794 0 471850 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 173346 0 173402 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 181994 0 182050 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 193586 0 193642 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 199382 0 199438 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 208122 0 208178 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 210974 0 211030 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 225510 0 225566 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 228362 0 228418 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 231306 0 231362 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 234158 0 234214 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 237102 0 237158 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 239954 0 240010 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 242898 0 242954 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 245750 0 245806 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 248694 0 248750 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 251546 0 251602 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 257342 0 257398 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 260286 0 260342 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 263138 0 263194 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 266082 0 266138 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 271878 0 271934 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 274730 0 274786 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 277674 0 277730 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 280526 0 280582 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 283470 0 283526 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 286322 0 286378 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 289266 0 289322 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 292118 0 292174 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 295062 0 295118 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 297914 0 297970 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 300858 0 300914 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 303710 0 303766 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 306654 0 306710 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 312450 0 312506 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 315302 0 315358 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 318246 0 318302 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 321098 0 321154 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 324042 0 324098 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 326894 0 326950 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 329838 0 329894 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 332690 0 332746 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 335634 0 335690 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 338486 0 338542 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 341430 0 341486 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 344282 0 344338 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 347226 0 347282 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 350078 0 350134 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 353022 0 353078 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 355874 0 355930 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 358818 0 358874 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 361670 0 361726 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 364614 0 364670 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 367466 0 367522 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 370410 0 370466 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 373262 0 373318 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 376206 0 376262 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 379058 0 379114 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 382002 0 382058 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 384854 0 384910 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 387798 0 387854 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 390650 0 390706 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 394514 0 394570 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 397458 0 397514 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 400310 0 400366 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 403254 0 403310 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 406106 0 406162 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 414846 0 414902 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 417698 0 417754 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 420642 0 420698 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 423494 0 423550 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 426438 0 426494 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 429290 0 429346 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 432234 0 432290 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 435086 0 435142 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 438030 0 438086 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 440882 0 440938 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 443826 0 443882 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 446678 0 446734 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 449622 0 449678 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 452474 0 452530 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 455418 0 455474 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 458270 0 458326 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 461214 0 461270 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 464066 0 464122 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 467010 0 467066 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 469862 0 469918 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 472806 0 472862 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 209042 0 209098 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 235170 0 235226 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 255410 0 255466 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 272798 0 272854 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 278594 0 278650 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 281538 0 281594 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 287334 0 287390 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 290186 0 290242 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 293130 0 293186 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 298926 0 298982 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 301778 0 301834 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 304722 0 304778 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 307574 0 307630 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 310518 0 310574 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 313370 0 313426 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 316314 0 316370 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 319166 0 319222 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 322110 0 322166 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 324962 0 325018 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 327906 0 327962 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 330758 0 330814 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 333702 0 333758 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 336554 0 336610 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 339498 0 339554 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 342350 0 342406 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 345294 0 345350 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 348146 0 348202 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 351090 0 351146 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 353942 0 353998 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 356886 0 356942 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 362682 0 362738 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 368478 0 368534 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 371330 0 371386 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 374274 0 374330 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 377126 0 377182 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 380070 0 380126 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 382922 0 382978 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 385866 0 385922 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 391662 0 391718 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 570704 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 570704 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 570704 6 vssd1
port 503 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 476207 573151
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 617058524
string GDS_START 1779578
<< end >>

