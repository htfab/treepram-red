magic
tech sky130A
magscale 1 2
timestamp 1636733283
<< obsli1 >>
rect 1104 2159 289955 290513
<< obsm1 >>
rect 290 1300 290614 290896
<< metal2 >>
rect 1214 292235 1270 293035
rect 3698 292235 3754 293035
rect 6274 292235 6330 293035
rect 8850 292235 8906 293035
rect 11334 292235 11390 293035
rect 13910 292235 13966 293035
rect 16486 292235 16542 293035
rect 19062 292235 19118 293035
rect 21546 292235 21602 293035
rect 24122 292235 24178 293035
rect 26698 292235 26754 293035
rect 29274 292235 29330 293035
rect 31758 292235 31814 293035
rect 34334 292235 34390 293035
rect 36910 292235 36966 293035
rect 39486 292235 39542 293035
rect 41970 292235 42026 293035
rect 44546 292235 44602 293035
rect 47122 292235 47178 293035
rect 49698 292235 49754 293035
rect 52182 292235 52238 293035
rect 54758 292235 54814 293035
rect 57334 292235 57390 293035
rect 59818 292235 59874 293035
rect 62394 292235 62450 293035
rect 64970 292235 65026 293035
rect 67546 292235 67602 293035
rect 70030 292235 70086 293035
rect 72606 292235 72662 293035
rect 75182 292235 75238 293035
rect 77758 292235 77814 293035
rect 80242 292235 80298 293035
rect 82818 292235 82874 293035
rect 85394 292235 85450 293035
rect 87970 292235 88026 293035
rect 90454 292235 90510 293035
rect 93030 292235 93086 293035
rect 95606 292235 95662 293035
rect 98182 292235 98238 293035
rect 100666 292235 100722 293035
rect 103242 292235 103298 293035
rect 105818 292235 105874 293035
rect 108302 292235 108358 293035
rect 110878 292235 110934 293035
rect 113454 292235 113510 293035
rect 116030 292235 116086 293035
rect 118514 292235 118570 293035
rect 121090 292235 121146 293035
rect 123666 292235 123722 293035
rect 126242 292235 126298 293035
rect 128726 292235 128782 293035
rect 131302 292235 131358 293035
rect 133878 292235 133934 293035
rect 136454 292235 136510 293035
rect 138938 292235 138994 293035
rect 141514 292235 141570 293035
rect 144090 292235 144146 293035
rect 146666 292235 146722 293035
rect 149150 292235 149206 293035
rect 151726 292235 151782 293035
rect 154302 292235 154358 293035
rect 156786 292235 156842 293035
rect 159362 292235 159418 293035
rect 161938 292235 161994 293035
rect 164514 292235 164570 293035
rect 166998 292235 167054 293035
rect 169574 292235 169630 293035
rect 172150 292235 172206 293035
rect 174726 292235 174782 293035
rect 177210 292235 177266 293035
rect 179786 292235 179842 293035
rect 182362 292235 182418 293035
rect 184938 292235 184994 293035
rect 187422 292235 187478 293035
rect 189998 292235 190054 293035
rect 192574 292235 192630 293035
rect 195150 292235 195206 293035
rect 197634 292235 197690 293035
rect 200210 292235 200266 293035
rect 202786 292235 202842 293035
rect 205270 292235 205326 293035
rect 207846 292235 207902 293035
rect 210422 292235 210478 293035
rect 212998 292235 213054 293035
rect 215482 292235 215538 293035
rect 218058 292235 218114 293035
rect 220634 292235 220690 293035
rect 223210 292235 223266 293035
rect 225694 292235 225750 293035
rect 228270 292235 228326 293035
rect 230846 292235 230902 293035
rect 233422 292235 233478 293035
rect 235906 292235 235962 293035
rect 238482 292235 238538 293035
rect 241058 292235 241114 293035
rect 243634 292235 243690 293035
rect 246118 292235 246174 293035
rect 248694 292235 248750 293035
rect 251270 292235 251326 293035
rect 253754 292235 253810 293035
rect 256330 292235 256386 293035
rect 258906 292235 258962 293035
rect 261482 292235 261538 293035
rect 263966 292235 264022 293035
rect 266542 292235 266598 293035
rect 269118 292235 269174 293035
rect 271694 292235 271750 293035
rect 274178 292235 274234 293035
rect 276754 292235 276810 293035
rect 279330 292235 279386 293035
rect 281906 292235 281962 293035
rect 284390 292235 284446 293035
rect 286966 292235 287022 293035
rect 289542 292235 289598 293035
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4986 0 5042 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 17958 0 18014 800
rect 18510 0 18566 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22098 0 22154 800
rect 22650 0 22706 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 25042 0 25098 800
rect 25594 0 25650 800
rect 26238 0 26294 800
rect 26790 0 26846 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30378 0 30434 800
rect 30930 0 30986 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34518 0 34574 800
rect 35070 0 35126 800
rect 35622 0 35678 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 40958 0 41014 800
rect 41510 0 41566 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43350 0 43406 800
rect 43902 0 43958 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46294 0 46350 800
rect 46846 0 46902 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56322 0 56378 800
rect 56874 0 56930 800
rect 57518 0 57574 800
rect 58070 0 58126 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59818 0 59874 800
rect 60462 0 60518 800
rect 61014 0 61070 800
rect 61658 0 61714 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64602 0 64658 800
rect 65154 0 65210 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66902 0 66958 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68742 0 68798 800
rect 69294 0 69350 800
rect 69846 0 69902 800
rect 70490 0 70546 800
rect 71042 0 71098 800
rect 71686 0 71742 800
rect 72238 0 72294 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75734 0 75790 800
rect 76378 0 76434 800
rect 76930 0 76986 800
rect 77574 0 77630 800
rect 78126 0 78182 800
rect 78770 0 78826 800
rect 79322 0 79378 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81070 0 81126 800
rect 81714 0 81770 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83462 0 83518 800
rect 84014 0 84070 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88154 0 88210 800
rect 88798 0 88854 800
rect 89350 0 89406 800
rect 89902 0 89958 800
rect 90546 0 90602 800
rect 91098 0 91154 800
rect 91742 0 91798 800
rect 92294 0 92350 800
rect 92846 0 92902 800
rect 93490 0 93546 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95238 0 95294 800
rect 95882 0 95938 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97630 0 97686 800
rect 98182 0 98238 800
rect 98826 0 98882 800
rect 99378 0 99434 800
rect 99930 0 99986 800
rect 100574 0 100630 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102322 0 102378 800
rect 102966 0 103022 800
rect 103518 0 103574 800
rect 104070 0 104126 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105910 0 105966 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107658 0 107714 800
rect 108210 0 108266 800
rect 108854 0 108910 800
rect 109406 0 109462 800
rect 109958 0 110014 800
rect 110602 0 110658 800
rect 111154 0 111210 800
rect 111798 0 111854 800
rect 112350 0 112406 800
rect 112994 0 113050 800
rect 113546 0 113602 800
rect 114098 0 114154 800
rect 114742 0 114798 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118882 0 118938 800
rect 119434 0 119490 800
rect 120078 0 120134 800
rect 120630 0 120686 800
rect 121182 0 121238 800
rect 121826 0 121882 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124770 0 124826 800
rect 125322 0 125378 800
rect 125966 0 126022 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127714 0 127770 800
rect 128266 0 128322 800
rect 128910 0 128966 800
rect 129462 0 129518 800
rect 130106 0 130162 800
rect 130658 0 130714 800
rect 131210 0 131266 800
rect 131854 0 131910 800
rect 132406 0 132462 800
rect 133050 0 133106 800
rect 133602 0 133658 800
rect 134154 0 134210 800
rect 134798 0 134854 800
rect 135350 0 135406 800
rect 135994 0 136050 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137742 0 137798 800
rect 138294 0 138350 800
rect 138938 0 138994 800
rect 139490 0 139546 800
rect 140134 0 140190 800
rect 140686 0 140742 800
rect 141238 0 141294 800
rect 141882 0 141938 800
rect 142434 0 142490 800
rect 143078 0 143134 800
rect 143630 0 143686 800
rect 144182 0 144238 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 146022 0 146078 800
rect 146574 0 146630 800
rect 147218 0 147274 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148966 0 149022 800
rect 149518 0 149574 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151266 0 151322 800
rect 151910 0 151966 800
rect 152462 0 152518 800
rect 153106 0 153162 800
rect 153658 0 153714 800
rect 154302 0 154358 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158350 0 158406 800
rect 158994 0 159050 800
rect 159546 0 159602 800
rect 160190 0 160246 800
rect 160742 0 160798 800
rect 161294 0 161350 800
rect 161938 0 161994 800
rect 162490 0 162546 800
rect 163134 0 163190 800
rect 163686 0 163742 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 166078 0 166134 800
rect 166630 0 166686 800
rect 167274 0 167330 800
rect 167826 0 167882 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169574 0 169630 800
rect 170218 0 170274 800
rect 170770 0 170826 800
rect 171414 0 171470 800
rect 171966 0 172022 800
rect 172518 0 172574 800
rect 173162 0 173218 800
rect 173714 0 173770 800
rect 174358 0 174414 800
rect 174910 0 174966 800
rect 175462 0 175518 800
rect 176106 0 176162 800
rect 176658 0 176714 800
rect 177302 0 177358 800
rect 177854 0 177910 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180246 0 180302 800
rect 180798 0 180854 800
rect 181442 0 181498 800
rect 181994 0 182050 800
rect 182546 0 182602 800
rect 183190 0 183246 800
rect 183742 0 183798 800
rect 184386 0 184442 800
rect 184938 0 184994 800
rect 185490 0 185546 800
rect 186134 0 186190 800
rect 186686 0 186742 800
rect 187330 0 187386 800
rect 187882 0 187938 800
rect 188526 0 188582 800
rect 189078 0 189134 800
rect 189630 0 189686 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191470 0 191526 800
rect 192022 0 192078 800
rect 192574 0 192630 800
rect 193218 0 193274 800
rect 193770 0 193826 800
rect 194414 0 194470 800
rect 194966 0 195022 800
rect 195518 0 195574 800
rect 196162 0 196218 800
rect 196714 0 196770 800
rect 197358 0 197414 800
rect 197910 0 197966 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201498 0 201554 800
rect 202050 0 202106 800
rect 202602 0 202658 800
rect 203246 0 203302 800
rect 203798 0 203854 800
rect 204442 0 204498 800
rect 204994 0 205050 800
rect 205638 0 205694 800
rect 206190 0 206246 800
rect 206742 0 206798 800
rect 207386 0 207442 800
rect 207938 0 207994 800
rect 208582 0 208638 800
rect 209134 0 209190 800
rect 209686 0 209742 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211526 0 211582 800
rect 212078 0 212134 800
rect 212630 0 212686 800
rect 213274 0 213330 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215022 0 215078 800
rect 215666 0 215722 800
rect 216218 0 216274 800
rect 216770 0 216826 800
rect 217414 0 217470 800
rect 217966 0 218022 800
rect 218610 0 218666 800
rect 219162 0 219218 800
rect 219714 0 219770 800
rect 220358 0 220414 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222750 0 222806 800
rect 223302 0 223358 800
rect 223854 0 223910 800
rect 224498 0 224554 800
rect 225050 0 225106 800
rect 225694 0 225750 800
rect 226246 0 226302 800
rect 226798 0 226854 800
rect 227442 0 227498 800
rect 227994 0 228050 800
rect 228638 0 228694 800
rect 229190 0 229246 800
rect 229742 0 229798 800
rect 230386 0 230442 800
rect 230938 0 230994 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234526 0 234582 800
rect 235078 0 235134 800
rect 235722 0 235778 800
rect 236274 0 236330 800
rect 236826 0 236882 800
rect 237470 0 237526 800
rect 238022 0 238078 800
rect 238666 0 238722 800
rect 239218 0 239274 800
rect 239862 0 239918 800
rect 240414 0 240470 800
rect 240966 0 241022 800
rect 241610 0 241666 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 243358 0 243414 800
rect 243910 0 243966 800
rect 244554 0 244610 800
rect 245106 0 245162 800
rect 245750 0 245806 800
rect 246302 0 246358 800
rect 246854 0 246910 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248694 0 248750 800
rect 249246 0 249302 800
rect 249890 0 249946 800
rect 250442 0 250498 800
rect 250994 0 251050 800
rect 251638 0 251694 800
rect 252190 0 252246 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 253938 0 253994 800
rect 254582 0 254638 800
rect 255134 0 255190 800
rect 255778 0 255834 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257526 0 257582 800
rect 258078 0 258134 800
rect 258722 0 258778 800
rect 259274 0 259330 800
rect 259918 0 259974 800
rect 260470 0 260526 800
rect 261022 0 261078 800
rect 261666 0 261722 800
rect 262218 0 262274 800
rect 262862 0 262918 800
rect 263414 0 263470 800
rect 263966 0 264022 800
rect 264610 0 264666 800
rect 265162 0 265218 800
rect 265806 0 265862 800
rect 266358 0 266414 800
rect 267002 0 267058 800
rect 267554 0 267610 800
rect 268106 0 268162 800
rect 268750 0 268806 800
rect 269302 0 269358 800
rect 269946 0 270002 800
rect 270498 0 270554 800
rect 271050 0 271106 800
rect 271694 0 271750 800
rect 272246 0 272302 800
rect 272890 0 272946 800
rect 273442 0 273498 800
rect 274086 0 274142 800
rect 274638 0 274694 800
rect 275190 0 275246 800
rect 275834 0 275890 800
rect 276386 0 276442 800
rect 277030 0 277086 800
rect 277582 0 277638 800
rect 278134 0 278190 800
rect 278778 0 278834 800
rect 279330 0 279386 800
rect 279974 0 280030 800
rect 280526 0 280582 800
rect 281078 0 281134 800
rect 281722 0 281778 800
rect 282274 0 282330 800
rect 282918 0 282974 800
rect 283470 0 283526 800
rect 284114 0 284170 800
rect 284666 0 284722 800
rect 285218 0 285274 800
rect 285862 0 285918 800
rect 286414 0 286470 800
rect 287058 0 287114 800
rect 287610 0 287666 800
rect 288162 0 288218 800
rect 288806 0 288862 800
rect 289358 0 289414 800
rect 290002 0 290058 800
rect 290554 0 290610 800
<< obsm2 >>
rect 296 292179 1158 292235
rect 1326 292179 3642 292235
rect 3810 292179 6218 292235
rect 6386 292179 8794 292235
rect 8962 292179 11278 292235
rect 11446 292179 13854 292235
rect 14022 292179 16430 292235
rect 16598 292179 19006 292235
rect 19174 292179 21490 292235
rect 21658 292179 24066 292235
rect 24234 292179 26642 292235
rect 26810 292179 29218 292235
rect 29386 292179 31702 292235
rect 31870 292179 34278 292235
rect 34446 292179 36854 292235
rect 37022 292179 39430 292235
rect 39598 292179 41914 292235
rect 42082 292179 44490 292235
rect 44658 292179 47066 292235
rect 47234 292179 49642 292235
rect 49810 292179 52126 292235
rect 52294 292179 54702 292235
rect 54870 292179 57278 292235
rect 57446 292179 59762 292235
rect 59930 292179 62338 292235
rect 62506 292179 64914 292235
rect 65082 292179 67490 292235
rect 67658 292179 69974 292235
rect 70142 292179 72550 292235
rect 72718 292179 75126 292235
rect 75294 292179 77702 292235
rect 77870 292179 80186 292235
rect 80354 292179 82762 292235
rect 82930 292179 85338 292235
rect 85506 292179 87914 292235
rect 88082 292179 90398 292235
rect 90566 292179 92974 292235
rect 93142 292179 95550 292235
rect 95718 292179 98126 292235
rect 98294 292179 100610 292235
rect 100778 292179 103186 292235
rect 103354 292179 105762 292235
rect 105930 292179 108246 292235
rect 108414 292179 110822 292235
rect 110990 292179 113398 292235
rect 113566 292179 115974 292235
rect 116142 292179 118458 292235
rect 118626 292179 121034 292235
rect 121202 292179 123610 292235
rect 123778 292179 126186 292235
rect 126354 292179 128670 292235
rect 128838 292179 131246 292235
rect 131414 292179 133822 292235
rect 133990 292179 136398 292235
rect 136566 292179 138882 292235
rect 139050 292179 141458 292235
rect 141626 292179 144034 292235
rect 144202 292179 146610 292235
rect 146778 292179 149094 292235
rect 149262 292179 151670 292235
rect 151838 292179 154246 292235
rect 154414 292179 156730 292235
rect 156898 292179 159306 292235
rect 159474 292179 161882 292235
rect 162050 292179 164458 292235
rect 164626 292179 166942 292235
rect 167110 292179 169518 292235
rect 169686 292179 172094 292235
rect 172262 292179 174670 292235
rect 174838 292179 177154 292235
rect 177322 292179 179730 292235
rect 179898 292179 182306 292235
rect 182474 292179 184882 292235
rect 185050 292179 187366 292235
rect 187534 292179 189942 292235
rect 190110 292179 192518 292235
rect 192686 292179 195094 292235
rect 195262 292179 197578 292235
rect 197746 292179 200154 292235
rect 200322 292179 202730 292235
rect 202898 292179 205214 292235
rect 205382 292179 207790 292235
rect 207958 292179 210366 292235
rect 210534 292179 212942 292235
rect 213110 292179 215426 292235
rect 215594 292179 218002 292235
rect 218170 292179 220578 292235
rect 220746 292179 223154 292235
rect 223322 292179 225638 292235
rect 225806 292179 228214 292235
rect 228382 292179 230790 292235
rect 230958 292179 233366 292235
rect 233534 292179 235850 292235
rect 236018 292179 238426 292235
rect 238594 292179 241002 292235
rect 241170 292179 243578 292235
rect 243746 292179 246062 292235
rect 246230 292179 248638 292235
rect 248806 292179 251214 292235
rect 251382 292179 253698 292235
rect 253866 292179 256274 292235
rect 256442 292179 258850 292235
rect 259018 292179 261426 292235
rect 261594 292179 263910 292235
rect 264078 292179 266486 292235
rect 266654 292179 269062 292235
rect 269230 292179 271638 292235
rect 271806 292179 274122 292235
rect 274290 292179 276698 292235
rect 276866 292179 279274 292235
rect 279442 292179 281850 292235
rect 282018 292179 284334 292235
rect 284502 292179 286910 292235
rect 287078 292179 289486 292235
rect 289654 292179 290608 292235
rect 296 856 290608 292179
rect 406 734 790 856
rect 958 734 1342 856
rect 1510 734 1986 856
rect 2154 734 2538 856
rect 2706 734 3182 856
rect 3350 734 3734 856
rect 3902 734 4286 856
rect 4454 734 4930 856
rect 5098 734 5482 856
rect 5650 734 6126 856
rect 6294 734 6678 856
rect 6846 734 7230 856
rect 7398 734 7874 856
rect 8042 734 8426 856
rect 8594 734 9070 856
rect 9238 734 9622 856
rect 9790 734 10266 856
rect 10434 734 10818 856
rect 10986 734 11370 856
rect 11538 734 12014 856
rect 12182 734 12566 856
rect 12734 734 13210 856
rect 13378 734 13762 856
rect 13930 734 14314 856
rect 14482 734 14958 856
rect 15126 734 15510 856
rect 15678 734 16154 856
rect 16322 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17902 856
rect 18070 734 18454 856
rect 18622 734 19098 856
rect 19266 734 19650 856
rect 19818 734 20294 856
rect 20462 734 20846 856
rect 21014 734 21398 856
rect 21566 734 22042 856
rect 22210 734 22594 856
rect 22762 734 23238 856
rect 23406 734 23790 856
rect 23958 734 24342 856
rect 24510 734 24986 856
rect 25154 734 25538 856
rect 25706 734 26182 856
rect 26350 734 26734 856
rect 26902 734 27378 856
rect 27546 734 27930 856
rect 28098 734 28482 856
rect 28650 734 29126 856
rect 29294 734 29678 856
rect 29846 734 30322 856
rect 30490 734 30874 856
rect 31042 734 31426 856
rect 31594 734 32070 856
rect 32238 734 32622 856
rect 32790 734 33266 856
rect 33434 734 33818 856
rect 33986 734 34462 856
rect 34630 734 35014 856
rect 35182 734 35566 856
rect 35734 734 36210 856
rect 36378 734 36762 856
rect 36930 734 37406 856
rect 37574 734 37958 856
rect 38126 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39706 856
rect 39874 734 40350 856
rect 40518 734 40902 856
rect 41070 734 41454 856
rect 41622 734 42098 856
rect 42266 734 42650 856
rect 42818 734 43294 856
rect 43462 734 43846 856
rect 44014 734 44490 856
rect 44658 734 45042 856
rect 45210 734 45594 856
rect 45762 734 46238 856
rect 46406 734 46790 856
rect 46958 734 47434 856
rect 47602 734 47986 856
rect 48154 734 48538 856
rect 48706 734 49182 856
rect 49350 734 49734 856
rect 49902 734 50378 856
rect 50546 734 50930 856
rect 51098 734 51574 856
rect 51742 734 52126 856
rect 52294 734 52678 856
rect 52846 734 53322 856
rect 53490 734 53874 856
rect 54042 734 54518 856
rect 54686 734 55070 856
rect 55238 734 55622 856
rect 55790 734 56266 856
rect 56434 734 56818 856
rect 56986 734 57462 856
rect 57630 734 58014 856
rect 58182 734 58566 856
rect 58734 734 59210 856
rect 59378 734 59762 856
rect 59930 734 60406 856
rect 60574 734 60958 856
rect 61126 734 61602 856
rect 61770 734 62154 856
rect 62322 734 62706 856
rect 62874 734 63350 856
rect 63518 734 63902 856
rect 64070 734 64546 856
rect 64714 734 65098 856
rect 65266 734 65650 856
rect 65818 734 66294 856
rect 66462 734 66846 856
rect 67014 734 67490 856
rect 67658 734 68042 856
rect 68210 734 68686 856
rect 68854 734 69238 856
rect 69406 734 69790 856
rect 69958 734 70434 856
rect 70602 734 70986 856
rect 71154 734 71630 856
rect 71798 734 72182 856
rect 72350 734 72734 856
rect 72902 734 73378 856
rect 73546 734 73930 856
rect 74098 734 74574 856
rect 74742 734 75126 856
rect 75294 734 75678 856
rect 75846 734 76322 856
rect 76490 734 76874 856
rect 77042 734 77518 856
rect 77686 734 78070 856
rect 78238 734 78714 856
rect 78882 734 79266 856
rect 79434 734 79818 856
rect 79986 734 80462 856
rect 80630 734 81014 856
rect 81182 734 81658 856
rect 81826 734 82210 856
rect 82378 734 82762 856
rect 82930 734 83406 856
rect 83574 734 83958 856
rect 84126 734 84602 856
rect 84770 734 85154 856
rect 85322 734 85798 856
rect 85966 734 86350 856
rect 86518 734 86902 856
rect 87070 734 87546 856
rect 87714 734 88098 856
rect 88266 734 88742 856
rect 88910 734 89294 856
rect 89462 734 89846 856
rect 90014 734 90490 856
rect 90658 734 91042 856
rect 91210 734 91686 856
rect 91854 734 92238 856
rect 92406 734 92790 856
rect 92958 734 93434 856
rect 93602 734 93986 856
rect 94154 734 94630 856
rect 94798 734 95182 856
rect 95350 734 95826 856
rect 95994 734 96378 856
rect 96546 734 96930 856
rect 97098 734 97574 856
rect 97742 734 98126 856
rect 98294 734 98770 856
rect 98938 734 99322 856
rect 99490 734 99874 856
rect 100042 734 100518 856
rect 100686 734 101070 856
rect 101238 734 101714 856
rect 101882 734 102266 856
rect 102434 734 102910 856
rect 103078 734 103462 856
rect 103630 734 104014 856
rect 104182 734 104658 856
rect 104826 734 105210 856
rect 105378 734 105854 856
rect 106022 734 106406 856
rect 106574 734 106958 856
rect 107126 734 107602 856
rect 107770 734 108154 856
rect 108322 734 108798 856
rect 108966 734 109350 856
rect 109518 734 109902 856
rect 110070 734 110546 856
rect 110714 734 111098 856
rect 111266 734 111742 856
rect 111910 734 112294 856
rect 112462 734 112938 856
rect 113106 734 113490 856
rect 113658 734 114042 856
rect 114210 734 114686 856
rect 114854 734 115238 856
rect 115406 734 115882 856
rect 116050 734 116434 856
rect 116602 734 116986 856
rect 117154 734 117630 856
rect 117798 734 118182 856
rect 118350 734 118826 856
rect 118994 734 119378 856
rect 119546 734 120022 856
rect 120190 734 120574 856
rect 120742 734 121126 856
rect 121294 734 121770 856
rect 121938 734 122322 856
rect 122490 734 122966 856
rect 123134 734 123518 856
rect 123686 734 124070 856
rect 124238 734 124714 856
rect 124882 734 125266 856
rect 125434 734 125910 856
rect 126078 734 126462 856
rect 126630 734 127014 856
rect 127182 734 127658 856
rect 127826 734 128210 856
rect 128378 734 128854 856
rect 129022 734 129406 856
rect 129574 734 130050 856
rect 130218 734 130602 856
rect 130770 734 131154 856
rect 131322 734 131798 856
rect 131966 734 132350 856
rect 132518 734 132994 856
rect 133162 734 133546 856
rect 133714 734 134098 856
rect 134266 734 134742 856
rect 134910 734 135294 856
rect 135462 734 135938 856
rect 136106 734 136490 856
rect 136658 734 137134 856
rect 137302 734 137686 856
rect 137854 734 138238 856
rect 138406 734 138882 856
rect 139050 734 139434 856
rect 139602 734 140078 856
rect 140246 734 140630 856
rect 140798 734 141182 856
rect 141350 734 141826 856
rect 141994 734 142378 856
rect 142546 734 143022 856
rect 143190 734 143574 856
rect 143742 734 144126 856
rect 144294 734 144770 856
rect 144938 734 145322 856
rect 145490 734 145966 856
rect 146134 734 146518 856
rect 146686 734 147162 856
rect 147330 734 147714 856
rect 147882 734 148266 856
rect 148434 734 148910 856
rect 149078 734 149462 856
rect 149630 734 150106 856
rect 150274 734 150658 856
rect 150826 734 151210 856
rect 151378 734 151854 856
rect 152022 734 152406 856
rect 152574 734 153050 856
rect 153218 734 153602 856
rect 153770 734 154246 856
rect 154414 734 154798 856
rect 154966 734 155350 856
rect 155518 734 155994 856
rect 156162 734 156546 856
rect 156714 734 157190 856
rect 157358 734 157742 856
rect 157910 734 158294 856
rect 158462 734 158938 856
rect 159106 734 159490 856
rect 159658 734 160134 856
rect 160302 734 160686 856
rect 160854 734 161238 856
rect 161406 734 161882 856
rect 162050 734 162434 856
rect 162602 734 163078 856
rect 163246 734 163630 856
rect 163798 734 164274 856
rect 164442 734 164826 856
rect 164994 734 165378 856
rect 165546 734 166022 856
rect 166190 734 166574 856
rect 166742 734 167218 856
rect 167386 734 167770 856
rect 167938 734 168322 856
rect 168490 734 168966 856
rect 169134 734 169518 856
rect 169686 734 170162 856
rect 170330 734 170714 856
rect 170882 734 171358 856
rect 171526 734 171910 856
rect 172078 734 172462 856
rect 172630 734 173106 856
rect 173274 734 173658 856
rect 173826 734 174302 856
rect 174470 734 174854 856
rect 175022 734 175406 856
rect 175574 734 176050 856
rect 176218 734 176602 856
rect 176770 734 177246 856
rect 177414 734 177798 856
rect 177966 734 178350 856
rect 178518 734 178994 856
rect 179162 734 179546 856
rect 179714 734 180190 856
rect 180358 734 180742 856
rect 180910 734 181386 856
rect 181554 734 181938 856
rect 182106 734 182490 856
rect 182658 734 183134 856
rect 183302 734 183686 856
rect 183854 734 184330 856
rect 184498 734 184882 856
rect 185050 734 185434 856
rect 185602 734 186078 856
rect 186246 734 186630 856
rect 186798 734 187274 856
rect 187442 734 187826 856
rect 187994 734 188470 856
rect 188638 734 189022 856
rect 189190 734 189574 856
rect 189742 734 190218 856
rect 190386 734 190770 856
rect 190938 734 191414 856
rect 191582 734 191966 856
rect 192134 734 192518 856
rect 192686 734 193162 856
rect 193330 734 193714 856
rect 193882 734 194358 856
rect 194526 734 194910 856
rect 195078 734 195462 856
rect 195630 734 196106 856
rect 196274 734 196658 856
rect 196826 734 197302 856
rect 197470 734 197854 856
rect 198022 734 198498 856
rect 198666 734 199050 856
rect 199218 734 199602 856
rect 199770 734 200246 856
rect 200414 734 200798 856
rect 200966 734 201442 856
rect 201610 734 201994 856
rect 202162 734 202546 856
rect 202714 734 203190 856
rect 203358 734 203742 856
rect 203910 734 204386 856
rect 204554 734 204938 856
rect 205106 734 205582 856
rect 205750 734 206134 856
rect 206302 734 206686 856
rect 206854 734 207330 856
rect 207498 734 207882 856
rect 208050 734 208526 856
rect 208694 734 209078 856
rect 209246 734 209630 856
rect 209798 734 210274 856
rect 210442 734 210826 856
rect 210994 734 211470 856
rect 211638 734 212022 856
rect 212190 734 212574 856
rect 212742 734 213218 856
rect 213386 734 213770 856
rect 213938 734 214414 856
rect 214582 734 214966 856
rect 215134 734 215610 856
rect 215778 734 216162 856
rect 216330 734 216714 856
rect 216882 734 217358 856
rect 217526 734 217910 856
rect 218078 734 218554 856
rect 218722 734 219106 856
rect 219274 734 219658 856
rect 219826 734 220302 856
rect 220470 734 220854 856
rect 221022 734 221498 856
rect 221666 734 222050 856
rect 222218 734 222694 856
rect 222862 734 223246 856
rect 223414 734 223798 856
rect 223966 734 224442 856
rect 224610 734 224994 856
rect 225162 734 225638 856
rect 225806 734 226190 856
rect 226358 734 226742 856
rect 226910 734 227386 856
rect 227554 734 227938 856
rect 228106 734 228582 856
rect 228750 734 229134 856
rect 229302 734 229686 856
rect 229854 734 230330 856
rect 230498 734 230882 856
rect 231050 734 231526 856
rect 231694 734 232078 856
rect 232246 734 232722 856
rect 232890 734 233274 856
rect 233442 734 233826 856
rect 233994 734 234470 856
rect 234638 734 235022 856
rect 235190 734 235666 856
rect 235834 734 236218 856
rect 236386 734 236770 856
rect 236938 734 237414 856
rect 237582 734 237966 856
rect 238134 734 238610 856
rect 238778 734 239162 856
rect 239330 734 239806 856
rect 239974 734 240358 856
rect 240526 734 240910 856
rect 241078 734 241554 856
rect 241722 734 242106 856
rect 242274 734 242750 856
rect 242918 734 243302 856
rect 243470 734 243854 856
rect 244022 734 244498 856
rect 244666 734 245050 856
rect 245218 734 245694 856
rect 245862 734 246246 856
rect 246414 734 246798 856
rect 246966 734 247442 856
rect 247610 734 247994 856
rect 248162 734 248638 856
rect 248806 734 249190 856
rect 249358 734 249834 856
rect 250002 734 250386 856
rect 250554 734 250938 856
rect 251106 734 251582 856
rect 251750 734 252134 856
rect 252302 734 252778 856
rect 252946 734 253330 856
rect 253498 734 253882 856
rect 254050 734 254526 856
rect 254694 734 255078 856
rect 255246 734 255722 856
rect 255890 734 256274 856
rect 256442 734 256918 856
rect 257086 734 257470 856
rect 257638 734 258022 856
rect 258190 734 258666 856
rect 258834 734 259218 856
rect 259386 734 259862 856
rect 260030 734 260414 856
rect 260582 734 260966 856
rect 261134 734 261610 856
rect 261778 734 262162 856
rect 262330 734 262806 856
rect 262974 734 263358 856
rect 263526 734 263910 856
rect 264078 734 264554 856
rect 264722 734 265106 856
rect 265274 734 265750 856
rect 265918 734 266302 856
rect 266470 734 266946 856
rect 267114 734 267498 856
rect 267666 734 268050 856
rect 268218 734 268694 856
rect 268862 734 269246 856
rect 269414 734 269890 856
rect 270058 734 270442 856
rect 270610 734 270994 856
rect 271162 734 271638 856
rect 271806 734 272190 856
rect 272358 734 272834 856
rect 273002 734 273386 856
rect 273554 734 274030 856
rect 274198 734 274582 856
rect 274750 734 275134 856
rect 275302 734 275778 856
rect 275946 734 276330 856
rect 276498 734 276974 856
rect 277142 734 277526 856
rect 277694 734 278078 856
rect 278246 734 278722 856
rect 278890 734 279274 856
rect 279442 734 279918 856
rect 280086 734 280470 856
rect 280638 734 281022 856
rect 281190 734 281666 856
rect 281834 734 282218 856
rect 282386 734 282862 856
rect 283030 734 283414 856
rect 283582 734 284058 856
rect 284226 734 284610 856
rect 284778 734 285162 856
rect 285330 734 285806 856
rect 285974 734 286358 856
rect 286526 734 287002 856
rect 287170 734 287554 856
rect 287722 734 288106 856
rect 288274 734 288750 856
rect 288918 734 289302 856
rect 289470 734 289946 856
rect 290114 734 290498 856
<< obsm3 >>
rect 1669 1395 288867 290529
<< metal4 >>
rect 4208 2128 4528 290544
rect 19568 2128 19888 290544
rect 34928 2128 35248 290544
rect 50288 2128 50608 290544
rect 65648 2128 65968 290544
rect 81008 2128 81328 290544
rect 96368 2128 96688 290544
rect 111728 2128 112048 290544
rect 127088 2128 127408 290544
rect 142448 2128 142768 290544
rect 157808 2128 158128 290544
rect 173168 2128 173488 290544
rect 188528 2128 188848 290544
rect 203888 2128 204208 290544
rect 219248 2128 219568 290544
rect 234608 2128 234928 290544
rect 249968 2128 250288 290544
rect 265328 2128 265648 290544
rect 280688 2128 281008 290544
<< obsm4 >>
rect 4659 3571 19488 290189
rect 19968 3571 34848 290189
rect 35328 3571 50208 290189
rect 50688 3571 65568 290189
rect 66048 3571 80928 290189
rect 81408 3571 96288 290189
rect 96768 3571 111648 290189
rect 112128 3571 127008 290189
rect 127488 3571 142368 290189
rect 142848 3571 157728 290189
rect 158208 3571 173088 290189
rect 173568 3571 188448 290189
rect 188928 3571 203808 290189
rect 204288 3571 219168 290189
rect 219648 3571 234528 290189
rect 235008 3571 249888 290189
rect 250368 3571 265248 290189
rect 265728 3571 280608 290189
rect 281088 3571 287901 290189
<< labels >>
rlabel metal2 s 1214 292235 1270 293035 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 77758 292235 77814 293035 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 85394 292235 85450 293035 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 93030 292235 93086 293035 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 100666 292235 100722 293035 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 108302 292235 108358 293035 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 116030 292235 116086 293035 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 123666 292235 123722 293035 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 131302 292235 131358 293035 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 138938 292235 138994 293035 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 146666 292235 146722 293035 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8850 292235 8906 293035 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 154302 292235 154358 293035 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 161938 292235 161994 293035 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 169574 292235 169630 293035 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 177210 292235 177266 293035 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 184938 292235 184994 293035 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 192574 292235 192630 293035 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 200210 292235 200266 293035 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 207846 292235 207902 293035 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 215482 292235 215538 293035 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 223210 292235 223266 293035 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 16486 292235 16542 293035 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 230846 292235 230902 293035 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 238482 292235 238538 293035 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 246118 292235 246174 293035 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 253754 292235 253810 293035 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 261482 292235 261538 293035 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 269118 292235 269174 293035 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 276754 292235 276810 293035 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 284390 292235 284446 293035 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24122 292235 24178 293035 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 31758 292235 31814 293035 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 39486 292235 39542 293035 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 47122 292235 47178 293035 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 54758 292235 54814 293035 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 62394 292235 62450 293035 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 70030 292235 70086 293035 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3698 292235 3754 293035 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 80242 292235 80298 293035 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 87970 292235 88026 293035 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 95606 292235 95662 293035 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 103242 292235 103298 293035 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 110878 292235 110934 293035 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 118514 292235 118570 293035 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 126242 292235 126298 293035 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 133878 292235 133934 293035 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 141514 292235 141570 293035 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 149150 292235 149206 293035 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11334 292235 11390 293035 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 156786 292235 156842 293035 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 164514 292235 164570 293035 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 172150 292235 172206 293035 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 179786 292235 179842 293035 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 187422 292235 187478 293035 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 195150 292235 195206 293035 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 202786 292235 202842 293035 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 210422 292235 210478 293035 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 218058 292235 218114 293035 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 225694 292235 225750 293035 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 19062 292235 19118 293035 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 233422 292235 233478 293035 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 241058 292235 241114 293035 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 248694 292235 248750 293035 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 256330 292235 256386 293035 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 263966 292235 264022 293035 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 271694 292235 271750 293035 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 279330 292235 279386 293035 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 286966 292235 287022 293035 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26698 292235 26754 293035 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 34334 292235 34390 293035 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 41970 292235 42026 293035 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 49698 292235 49754 293035 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 57334 292235 57390 293035 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 64970 292235 65026 293035 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 72606 292235 72662 293035 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6274 292235 6330 293035 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 82818 292235 82874 293035 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 90454 292235 90510 293035 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 98182 292235 98238 293035 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 105818 292235 105874 293035 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 113454 292235 113510 293035 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 121090 292235 121146 293035 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 128726 292235 128782 293035 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 136454 292235 136510 293035 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 144090 292235 144146 293035 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 151726 292235 151782 293035 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 13910 292235 13966 293035 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 159362 292235 159418 293035 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 166998 292235 167054 293035 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 174726 292235 174782 293035 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 182362 292235 182418 293035 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 189998 292235 190054 293035 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 197634 292235 197690 293035 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 205270 292235 205326 293035 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 212998 292235 213054 293035 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 220634 292235 220690 293035 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 228270 292235 228326 293035 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 21546 292235 21602 293035 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 235906 292235 235962 293035 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 243634 292235 243690 293035 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 251270 292235 251326 293035 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 258906 292235 258962 293035 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 266542 292235 266598 293035 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 274178 292235 274234 293035 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 281906 292235 281962 293035 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 289542 292235 289598 293035 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 29274 292235 29330 293035 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 36910 292235 36966 293035 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 44546 292235 44602 293035 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 52182 292235 52238 293035 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 59818 292235 59874 293035 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 67546 292235 67602 293035 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 75182 292235 75238 293035 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 289358 0 289414 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 290002 0 290058 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 290554 0 290610 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 248694 0 248750 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 255778 0 255834 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 262862 0 262918 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 275190 0 275246 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 280526 0 280582 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 282274 0 282330 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 285862 0 285918 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 240414 0 240470 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 243910 0 243966 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 245750 0 245806 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 247498 0 247554 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 249246 0 249302 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 250994 0 251050 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 254582 0 254638 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 258078 0 258134 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 261666 0 261722 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 263414 0 263470 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 265162 0 265218 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 267002 0 267058 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 268750 0 268806 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 270498 0 270554 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 272246 0 272302 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 274086 0 274142 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 275834 0 275890 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 277582 0 277638 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 279330 0 279386 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 281078 0 281134 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 282918 0 282974 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 284666 0 284722 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 286414 0 286470 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 288162 0 288218 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 158994 0 159050 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 171414 0 171470 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 176658 0 176714 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 181994 0 182050 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 183742 0 183798 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 187330 0 187386 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 204994 0 205050 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 208582 0 208638 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 210330 0 210386 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 212078 0 212134 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 217414 0 217470 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 224498 0 224554 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 226246 0 226302 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 229742 0 229798 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 236826 0 236882 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 238666 0 238722 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 242806 0 242862 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 244554 0 244610 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 263966 0 264022 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 265806 0 265862 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 269302 0 269358 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 278134 0 278190 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 281722 0 281778 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 288806 0 288862 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 230386 0 230442 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 239218 0 239274 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 290544 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 290544 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 290544 6 vssd1
port 503 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 290891 293035
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 218664374
string GDS_START 1742490
<< end >>

