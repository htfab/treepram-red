magic
tech sky130A
magscale 1 2
timestamp 1636730130
<< obsli1 >>
rect 1104 1377 199335 199665
<< obsm1 >>
rect 198 76 199626 200116
<< metal2 >>
rect 846 201156 902 201956
rect 2594 201156 2650 201956
rect 4342 201156 4398 201956
rect 6090 201156 6146 201956
rect 7838 201156 7894 201956
rect 9586 201156 9642 201956
rect 11334 201156 11390 201956
rect 13082 201156 13138 201956
rect 14830 201156 14886 201956
rect 16578 201156 16634 201956
rect 18326 201156 18382 201956
rect 20074 201156 20130 201956
rect 21822 201156 21878 201956
rect 23570 201156 23626 201956
rect 25318 201156 25374 201956
rect 27066 201156 27122 201956
rect 28814 201156 28870 201956
rect 30562 201156 30618 201956
rect 32310 201156 32366 201956
rect 34150 201156 34206 201956
rect 35898 201156 35954 201956
rect 37646 201156 37702 201956
rect 39394 201156 39450 201956
rect 41142 201156 41198 201956
rect 42890 201156 42946 201956
rect 44638 201156 44694 201956
rect 46386 201156 46442 201956
rect 48134 201156 48190 201956
rect 49882 201156 49938 201956
rect 51630 201156 51686 201956
rect 53378 201156 53434 201956
rect 55126 201156 55182 201956
rect 56874 201156 56930 201956
rect 58622 201156 58678 201956
rect 60370 201156 60426 201956
rect 62118 201156 62174 201956
rect 63866 201156 63922 201956
rect 65614 201156 65670 201956
rect 67454 201156 67510 201956
rect 69202 201156 69258 201956
rect 70950 201156 71006 201956
rect 72698 201156 72754 201956
rect 74446 201156 74502 201956
rect 76194 201156 76250 201956
rect 77942 201156 77998 201956
rect 79690 201156 79746 201956
rect 81438 201156 81494 201956
rect 83186 201156 83242 201956
rect 84934 201156 84990 201956
rect 86682 201156 86738 201956
rect 88430 201156 88486 201956
rect 90178 201156 90234 201956
rect 91926 201156 91982 201956
rect 93674 201156 93730 201956
rect 95422 201156 95478 201956
rect 97170 201156 97226 201956
rect 98918 201156 98974 201956
rect 100758 201156 100814 201956
rect 102506 201156 102562 201956
rect 104254 201156 104310 201956
rect 106002 201156 106058 201956
rect 107750 201156 107806 201956
rect 109498 201156 109554 201956
rect 111246 201156 111302 201956
rect 112994 201156 113050 201956
rect 114742 201156 114798 201956
rect 116490 201156 116546 201956
rect 118238 201156 118294 201956
rect 119986 201156 120042 201956
rect 121734 201156 121790 201956
rect 123482 201156 123538 201956
rect 125230 201156 125286 201956
rect 126978 201156 127034 201956
rect 128726 201156 128782 201956
rect 130474 201156 130530 201956
rect 132222 201156 132278 201956
rect 134062 201156 134118 201956
rect 135810 201156 135866 201956
rect 137558 201156 137614 201956
rect 139306 201156 139362 201956
rect 141054 201156 141110 201956
rect 142802 201156 142858 201956
rect 144550 201156 144606 201956
rect 146298 201156 146354 201956
rect 148046 201156 148102 201956
rect 149794 201156 149850 201956
rect 151542 201156 151598 201956
rect 153290 201156 153346 201956
rect 155038 201156 155094 201956
rect 156786 201156 156842 201956
rect 158534 201156 158590 201956
rect 160282 201156 160338 201956
rect 162030 201156 162086 201956
rect 163778 201156 163834 201956
rect 165526 201156 165582 201956
rect 167366 201156 167422 201956
rect 169114 201156 169170 201956
rect 170862 201156 170918 201956
rect 172610 201156 172666 201956
rect 174358 201156 174414 201956
rect 176106 201156 176162 201956
rect 177854 201156 177910 201956
rect 179602 201156 179658 201956
rect 181350 201156 181406 201956
rect 183098 201156 183154 201956
rect 184846 201156 184902 201956
rect 186594 201156 186650 201956
rect 188342 201156 188398 201956
rect 190090 201156 190146 201956
rect 191838 201156 191894 201956
rect 193586 201156 193642 201956
rect 195334 201156 195390 201956
rect 197082 201156 197138 201956
rect 198830 201156 198886 201956
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39486 0 39542 800
rect 39854 0 39910 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 62946 0 63002 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66994 0 67050 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88890 0 88946 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90178 0 90234 800
rect 90546 0 90602 800
rect 90914 0 90970 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121366 0 121422 800
rect 121734 0 121790 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130290 0 130346 800
rect 130658 0 130714 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142434 0 142490 800
rect 142802 0 142858 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155406 0 155462 800
rect 155774 0 155830 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158258 0 158314 800
rect 158626 0 158682 800
rect 159086 0 159142 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161110 0 161166 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 163134 0 163190 800
rect 163502 0 163558 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171230 0 171286 800
rect 171598 0 171654 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 174082 0 174138 800
rect 174450 0 174506 800
rect 174818 0 174874 800
rect 175278 0 175334 800
rect 175646 0 175702 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177302 0 177358 800
rect 177670 0 177726 800
rect 178130 0 178186 800
rect 178498 0 178554 800
rect 178866 0 178922 800
rect 179326 0 179382 800
rect 179694 0 179750 800
rect 180154 0 180210 800
rect 180522 0 180578 800
rect 180890 0 180946 800
rect 181350 0 181406 800
rect 181718 0 181774 800
rect 182178 0 182234 800
rect 182546 0 182602 800
rect 182914 0 182970 800
rect 183374 0 183430 800
rect 183742 0 183798 800
rect 184202 0 184258 800
rect 184570 0 184626 800
rect 184938 0 184994 800
rect 185398 0 185454 800
rect 185766 0 185822 800
rect 186226 0 186282 800
rect 186594 0 186650 800
rect 187054 0 187110 800
rect 187422 0 187478 800
rect 187790 0 187846 800
rect 188250 0 188306 800
rect 188618 0 188674 800
rect 189078 0 189134 800
rect 189446 0 189502 800
rect 189814 0 189870 800
rect 190274 0 190330 800
rect 190642 0 190698 800
rect 191102 0 191158 800
rect 191470 0 191526 800
rect 191838 0 191894 800
rect 192298 0 192354 800
rect 192666 0 192722 800
rect 193126 0 193182 800
rect 193494 0 193550 800
rect 193862 0 193918 800
rect 194322 0 194378 800
rect 194690 0 194746 800
rect 195150 0 195206 800
rect 195518 0 195574 800
rect 195886 0 195942 800
rect 196346 0 196402 800
rect 196714 0 196770 800
rect 197174 0 197230 800
rect 197542 0 197598 800
rect 197910 0 197966 800
rect 198370 0 198426 800
rect 198738 0 198794 800
rect 199198 0 199254 800
rect 199566 0 199622 800
<< obsm2 >>
rect 204 201100 790 201226
rect 958 201100 2538 201226
rect 2706 201100 4286 201226
rect 4454 201100 6034 201226
rect 6202 201100 7782 201226
rect 7950 201100 9530 201226
rect 9698 201100 11278 201226
rect 11446 201100 13026 201226
rect 13194 201100 14774 201226
rect 14942 201100 16522 201226
rect 16690 201100 18270 201226
rect 18438 201100 20018 201226
rect 20186 201100 21766 201226
rect 21934 201100 23514 201226
rect 23682 201100 25262 201226
rect 25430 201100 27010 201226
rect 27178 201100 28758 201226
rect 28926 201100 30506 201226
rect 30674 201100 32254 201226
rect 32422 201100 34094 201226
rect 34262 201100 35842 201226
rect 36010 201100 37590 201226
rect 37758 201100 39338 201226
rect 39506 201100 41086 201226
rect 41254 201100 42834 201226
rect 43002 201100 44582 201226
rect 44750 201100 46330 201226
rect 46498 201100 48078 201226
rect 48246 201100 49826 201226
rect 49994 201100 51574 201226
rect 51742 201100 53322 201226
rect 53490 201100 55070 201226
rect 55238 201100 56818 201226
rect 56986 201100 58566 201226
rect 58734 201100 60314 201226
rect 60482 201100 62062 201226
rect 62230 201100 63810 201226
rect 63978 201100 65558 201226
rect 65726 201100 67398 201226
rect 67566 201100 69146 201226
rect 69314 201100 70894 201226
rect 71062 201100 72642 201226
rect 72810 201100 74390 201226
rect 74558 201100 76138 201226
rect 76306 201100 77886 201226
rect 78054 201100 79634 201226
rect 79802 201100 81382 201226
rect 81550 201100 83130 201226
rect 83298 201100 84878 201226
rect 85046 201100 86626 201226
rect 86794 201100 88374 201226
rect 88542 201100 90122 201226
rect 90290 201100 91870 201226
rect 92038 201100 93618 201226
rect 93786 201100 95366 201226
rect 95534 201100 97114 201226
rect 97282 201100 98862 201226
rect 99030 201100 100702 201226
rect 100870 201100 102450 201226
rect 102618 201100 104198 201226
rect 104366 201100 105946 201226
rect 106114 201100 107694 201226
rect 107862 201100 109442 201226
rect 109610 201100 111190 201226
rect 111358 201100 112938 201226
rect 113106 201100 114686 201226
rect 114854 201100 116434 201226
rect 116602 201100 118182 201226
rect 118350 201100 119930 201226
rect 120098 201100 121678 201226
rect 121846 201100 123426 201226
rect 123594 201100 125174 201226
rect 125342 201100 126922 201226
rect 127090 201100 128670 201226
rect 128838 201100 130418 201226
rect 130586 201100 132166 201226
rect 132334 201100 134006 201226
rect 134174 201100 135754 201226
rect 135922 201100 137502 201226
rect 137670 201100 139250 201226
rect 139418 201100 140998 201226
rect 141166 201100 142746 201226
rect 142914 201100 144494 201226
rect 144662 201100 146242 201226
rect 146410 201100 147990 201226
rect 148158 201100 149738 201226
rect 149906 201100 151486 201226
rect 151654 201100 153234 201226
rect 153402 201100 154982 201226
rect 155150 201100 156730 201226
rect 156898 201100 158478 201226
rect 158646 201100 160226 201226
rect 160394 201100 161974 201226
rect 162142 201100 163722 201226
rect 163890 201100 165470 201226
rect 165638 201100 167310 201226
rect 167478 201100 169058 201226
rect 169226 201100 170806 201226
rect 170974 201100 172554 201226
rect 172722 201100 174302 201226
rect 174470 201100 176050 201226
rect 176218 201100 177798 201226
rect 177966 201100 179546 201226
rect 179714 201100 181294 201226
rect 181462 201100 183042 201226
rect 183210 201100 184790 201226
rect 184958 201100 186538 201226
rect 186706 201100 188286 201226
rect 188454 201100 190034 201226
rect 190202 201100 191782 201226
rect 191950 201100 193530 201226
rect 193698 201100 195278 201226
rect 195446 201100 197026 201226
rect 197194 201100 198774 201226
rect 198942 201100 199620 201226
rect 204 856 199620 201100
rect 314 70 514 856
rect 682 70 882 856
rect 1050 70 1342 856
rect 1510 70 1710 856
rect 1878 70 2170 856
rect 2338 70 2538 856
rect 2706 70 2906 856
rect 3074 70 3366 856
rect 3534 70 3734 856
rect 3902 70 4194 856
rect 4362 70 4562 856
rect 4730 70 4930 856
rect 5098 70 5390 856
rect 5558 70 5758 856
rect 5926 70 6218 856
rect 6386 70 6586 856
rect 6754 70 6954 856
rect 7122 70 7414 856
rect 7582 70 7782 856
rect 7950 70 8242 856
rect 8410 70 8610 856
rect 8778 70 8978 856
rect 9146 70 9438 856
rect 9606 70 9806 856
rect 9974 70 10266 856
rect 10434 70 10634 856
rect 10802 70 11002 856
rect 11170 70 11462 856
rect 11630 70 11830 856
rect 11998 70 12290 856
rect 12458 70 12658 856
rect 12826 70 13026 856
rect 13194 70 13486 856
rect 13654 70 13854 856
rect 14022 70 14314 856
rect 14482 70 14682 856
rect 14850 70 15142 856
rect 15310 70 15510 856
rect 15678 70 15878 856
rect 16046 70 16338 856
rect 16506 70 16706 856
rect 16874 70 17166 856
rect 17334 70 17534 856
rect 17702 70 17902 856
rect 18070 70 18362 856
rect 18530 70 18730 856
rect 18898 70 19190 856
rect 19358 70 19558 856
rect 19726 70 19926 856
rect 20094 70 20386 856
rect 20554 70 20754 856
rect 20922 70 21214 856
rect 21382 70 21582 856
rect 21750 70 21950 856
rect 22118 70 22410 856
rect 22578 70 22778 856
rect 22946 70 23238 856
rect 23406 70 23606 856
rect 23774 70 23974 856
rect 24142 70 24434 856
rect 24602 70 24802 856
rect 24970 70 25262 856
rect 25430 70 25630 856
rect 25798 70 25998 856
rect 26166 70 26458 856
rect 26626 70 26826 856
rect 26994 70 27286 856
rect 27454 70 27654 856
rect 27822 70 28022 856
rect 28190 70 28482 856
rect 28650 70 28850 856
rect 29018 70 29310 856
rect 29478 70 29678 856
rect 29846 70 30138 856
rect 30306 70 30506 856
rect 30674 70 30874 856
rect 31042 70 31334 856
rect 31502 70 31702 856
rect 31870 70 32162 856
rect 32330 70 32530 856
rect 32698 70 32898 856
rect 33066 70 33358 856
rect 33526 70 33726 856
rect 33894 70 34186 856
rect 34354 70 34554 856
rect 34722 70 34922 856
rect 35090 70 35382 856
rect 35550 70 35750 856
rect 35918 70 36210 856
rect 36378 70 36578 856
rect 36746 70 36946 856
rect 37114 70 37406 856
rect 37574 70 37774 856
rect 37942 70 38234 856
rect 38402 70 38602 856
rect 38770 70 38970 856
rect 39138 70 39430 856
rect 39598 70 39798 856
rect 39966 70 40258 856
rect 40426 70 40626 856
rect 40794 70 40994 856
rect 41162 70 41454 856
rect 41622 70 41822 856
rect 41990 70 42282 856
rect 42450 70 42650 856
rect 42818 70 43110 856
rect 43278 70 43478 856
rect 43646 70 43846 856
rect 44014 70 44306 856
rect 44474 70 44674 856
rect 44842 70 45134 856
rect 45302 70 45502 856
rect 45670 70 45870 856
rect 46038 70 46330 856
rect 46498 70 46698 856
rect 46866 70 47158 856
rect 47326 70 47526 856
rect 47694 70 47894 856
rect 48062 70 48354 856
rect 48522 70 48722 856
rect 48890 70 49182 856
rect 49350 70 49550 856
rect 49718 70 49918 856
rect 50086 70 50378 856
rect 50546 70 50746 856
rect 50914 70 51206 856
rect 51374 70 51574 856
rect 51742 70 51942 856
rect 52110 70 52402 856
rect 52570 70 52770 856
rect 52938 70 53230 856
rect 53398 70 53598 856
rect 53766 70 53966 856
rect 54134 70 54426 856
rect 54594 70 54794 856
rect 54962 70 55254 856
rect 55422 70 55622 856
rect 55790 70 55990 856
rect 56158 70 56450 856
rect 56618 70 56818 856
rect 56986 70 57278 856
rect 57446 70 57646 856
rect 57814 70 58106 856
rect 58274 70 58474 856
rect 58642 70 58842 856
rect 59010 70 59302 856
rect 59470 70 59670 856
rect 59838 70 60130 856
rect 60298 70 60498 856
rect 60666 70 60866 856
rect 61034 70 61326 856
rect 61494 70 61694 856
rect 61862 70 62154 856
rect 62322 70 62522 856
rect 62690 70 62890 856
rect 63058 70 63350 856
rect 63518 70 63718 856
rect 63886 70 64178 856
rect 64346 70 64546 856
rect 64714 70 64914 856
rect 65082 70 65374 856
rect 65542 70 65742 856
rect 65910 70 66202 856
rect 66370 70 66570 856
rect 66738 70 66938 856
rect 67106 70 67398 856
rect 67566 70 67766 856
rect 67934 70 68226 856
rect 68394 70 68594 856
rect 68762 70 68962 856
rect 69130 70 69422 856
rect 69590 70 69790 856
rect 69958 70 70250 856
rect 70418 70 70618 856
rect 70786 70 70986 856
rect 71154 70 71446 856
rect 71614 70 71814 856
rect 71982 70 72274 856
rect 72442 70 72642 856
rect 72810 70 73102 856
rect 73270 70 73470 856
rect 73638 70 73838 856
rect 74006 70 74298 856
rect 74466 70 74666 856
rect 74834 70 75126 856
rect 75294 70 75494 856
rect 75662 70 75862 856
rect 76030 70 76322 856
rect 76490 70 76690 856
rect 76858 70 77150 856
rect 77318 70 77518 856
rect 77686 70 77886 856
rect 78054 70 78346 856
rect 78514 70 78714 856
rect 78882 70 79174 856
rect 79342 70 79542 856
rect 79710 70 79910 856
rect 80078 70 80370 856
rect 80538 70 80738 856
rect 80906 70 81198 856
rect 81366 70 81566 856
rect 81734 70 81934 856
rect 82102 70 82394 856
rect 82562 70 82762 856
rect 82930 70 83222 856
rect 83390 70 83590 856
rect 83758 70 83958 856
rect 84126 70 84418 856
rect 84586 70 84786 856
rect 84954 70 85246 856
rect 85414 70 85614 856
rect 85782 70 86074 856
rect 86242 70 86442 856
rect 86610 70 86810 856
rect 86978 70 87270 856
rect 87438 70 87638 856
rect 87806 70 88098 856
rect 88266 70 88466 856
rect 88634 70 88834 856
rect 89002 70 89294 856
rect 89462 70 89662 856
rect 89830 70 90122 856
rect 90290 70 90490 856
rect 90658 70 90858 856
rect 91026 70 91318 856
rect 91486 70 91686 856
rect 91854 70 92146 856
rect 92314 70 92514 856
rect 92682 70 92882 856
rect 93050 70 93342 856
rect 93510 70 93710 856
rect 93878 70 94170 856
rect 94338 70 94538 856
rect 94706 70 94906 856
rect 95074 70 95366 856
rect 95534 70 95734 856
rect 95902 70 96194 856
rect 96362 70 96562 856
rect 96730 70 96930 856
rect 97098 70 97390 856
rect 97558 70 97758 856
rect 97926 70 98218 856
rect 98386 70 98586 856
rect 98754 70 98954 856
rect 99122 70 99414 856
rect 99582 70 99782 856
rect 99950 70 100242 856
rect 100410 70 100610 856
rect 100778 70 101070 856
rect 101238 70 101438 856
rect 101606 70 101806 856
rect 101974 70 102266 856
rect 102434 70 102634 856
rect 102802 70 103094 856
rect 103262 70 103462 856
rect 103630 70 103830 856
rect 103998 70 104290 856
rect 104458 70 104658 856
rect 104826 70 105118 856
rect 105286 70 105486 856
rect 105654 70 105854 856
rect 106022 70 106314 856
rect 106482 70 106682 856
rect 106850 70 107142 856
rect 107310 70 107510 856
rect 107678 70 107878 856
rect 108046 70 108338 856
rect 108506 70 108706 856
rect 108874 70 109166 856
rect 109334 70 109534 856
rect 109702 70 109902 856
rect 110070 70 110362 856
rect 110530 70 110730 856
rect 110898 70 111190 856
rect 111358 70 111558 856
rect 111726 70 111926 856
rect 112094 70 112386 856
rect 112554 70 112754 856
rect 112922 70 113214 856
rect 113382 70 113582 856
rect 113750 70 113950 856
rect 114118 70 114410 856
rect 114578 70 114778 856
rect 114946 70 115238 856
rect 115406 70 115606 856
rect 115774 70 116066 856
rect 116234 70 116434 856
rect 116602 70 116802 856
rect 116970 70 117262 856
rect 117430 70 117630 856
rect 117798 70 118090 856
rect 118258 70 118458 856
rect 118626 70 118826 856
rect 118994 70 119286 856
rect 119454 70 119654 856
rect 119822 70 120114 856
rect 120282 70 120482 856
rect 120650 70 120850 856
rect 121018 70 121310 856
rect 121478 70 121678 856
rect 121846 70 122138 856
rect 122306 70 122506 856
rect 122674 70 122874 856
rect 123042 70 123334 856
rect 123502 70 123702 856
rect 123870 70 124162 856
rect 124330 70 124530 856
rect 124698 70 124898 856
rect 125066 70 125358 856
rect 125526 70 125726 856
rect 125894 70 126186 856
rect 126354 70 126554 856
rect 126722 70 126922 856
rect 127090 70 127382 856
rect 127550 70 127750 856
rect 127918 70 128210 856
rect 128378 70 128578 856
rect 128746 70 129038 856
rect 129206 70 129406 856
rect 129574 70 129774 856
rect 129942 70 130234 856
rect 130402 70 130602 856
rect 130770 70 131062 856
rect 131230 70 131430 856
rect 131598 70 131798 856
rect 131966 70 132258 856
rect 132426 70 132626 856
rect 132794 70 133086 856
rect 133254 70 133454 856
rect 133622 70 133822 856
rect 133990 70 134282 856
rect 134450 70 134650 856
rect 134818 70 135110 856
rect 135278 70 135478 856
rect 135646 70 135846 856
rect 136014 70 136306 856
rect 136474 70 136674 856
rect 136842 70 137134 856
rect 137302 70 137502 856
rect 137670 70 137870 856
rect 138038 70 138330 856
rect 138498 70 138698 856
rect 138866 70 139158 856
rect 139326 70 139526 856
rect 139694 70 139894 856
rect 140062 70 140354 856
rect 140522 70 140722 856
rect 140890 70 141182 856
rect 141350 70 141550 856
rect 141718 70 141918 856
rect 142086 70 142378 856
rect 142546 70 142746 856
rect 142914 70 143206 856
rect 143374 70 143574 856
rect 143742 70 144034 856
rect 144202 70 144402 856
rect 144570 70 144770 856
rect 144938 70 145230 856
rect 145398 70 145598 856
rect 145766 70 146058 856
rect 146226 70 146426 856
rect 146594 70 146794 856
rect 146962 70 147254 856
rect 147422 70 147622 856
rect 147790 70 148082 856
rect 148250 70 148450 856
rect 148618 70 148818 856
rect 148986 70 149278 856
rect 149446 70 149646 856
rect 149814 70 150106 856
rect 150274 70 150474 856
rect 150642 70 150842 856
rect 151010 70 151302 856
rect 151470 70 151670 856
rect 151838 70 152130 856
rect 152298 70 152498 856
rect 152666 70 152866 856
rect 153034 70 153326 856
rect 153494 70 153694 856
rect 153862 70 154154 856
rect 154322 70 154522 856
rect 154690 70 154890 856
rect 155058 70 155350 856
rect 155518 70 155718 856
rect 155886 70 156178 856
rect 156346 70 156546 856
rect 156714 70 156914 856
rect 157082 70 157374 856
rect 157542 70 157742 856
rect 157910 70 158202 856
rect 158370 70 158570 856
rect 158738 70 159030 856
rect 159198 70 159398 856
rect 159566 70 159766 856
rect 159934 70 160226 856
rect 160394 70 160594 856
rect 160762 70 161054 856
rect 161222 70 161422 856
rect 161590 70 161790 856
rect 161958 70 162250 856
rect 162418 70 162618 856
rect 162786 70 163078 856
rect 163246 70 163446 856
rect 163614 70 163814 856
rect 163982 70 164274 856
rect 164442 70 164642 856
rect 164810 70 165102 856
rect 165270 70 165470 856
rect 165638 70 165838 856
rect 166006 70 166298 856
rect 166466 70 166666 856
rect 166834 70 167126 856
rect 167294 70 167494 856
rect 167662 70 167862 856
rect 168030 70 168322 856
rect 168490 70 168690 856
rect 168858 70 169150 856
rect 169318 70 169518 856
rect 169686 70 169886 856
rect 170054 70 170346 856
rect 170514 70 170714 856
rect 170882 70 171174 856
rect 171342 70 171542 856
rect 171710 70 172002 856
rect 172170 70 172370 856
rect 172538 70 172738 856
rect 172906 70 173198 856
rect 173366 70 173566 856
rect 173734 70 174026 856
rect 174194 70 174394 856
rect 174562 70 174762 856
rect 174930 70 175222 856
rect 175390 70 175590 856
rect 175758 70 176050 856
rect 176218 70 176418 856
rect 176586 70 176786 856
rect 176954 70 177246 856
rect 177414 70 177614 856
rect 177782 70 178074 856
rect 178242 70 178442 856
rect 178610 70 178810 856
rect 178978 70 179270 856
rect 179438 70 179638 856
rect 179806 70 180098 856
rect 180266 70 180466 856
rect 180634 70 180834 856
rect 181002 70 181294 856
rect 181462 70 181662 856
rect 181830 70 182122 856
rect 182290 70 182490 856
rect 182658 70 182858 856
rect 183026 70 183318 856
rect 183486 70 183686 856
rect 183854 70 184146 856
rect 184314 70 184514 856
rect 184682 70 184882 856
rect 185050 70 185342 856
rect 185510 70 185710 856
rect 185878 70 186170 856
rect 186338 70 186538 856
rect 186706 70 186998 856
rect 187166 70 187366 856
rect 187534 70 187734 856
rect 187902 70 188194 856
rect 188362 70 188562 856
rect 188730 70 189022 856
rect 189190 70 189390 856
rect 189558 70 189758 856
rect 189926 70 190218 856
rect 190386 70 190586 856
rect 190754 70 191046 856
rect 191214 70 191414 856
rect 191582 70 191782 856
rect 191950 70 192242 856
rect 192410 70 192610 856
rect 192778 70 193070 856
rect 193238 70 193438 856
rect 193606 70 193806 856
rect 193974 70 194266 856
rect 194434 70 194634 856
rect 194802 70 195094 856
rect 195262 70 195462 856
rect 195630 70 195830 856
rect 195998 70 196290 856
rect 196458 70 196658 856
rect 196826 70 197118 856
rect 197286 70 197486 856
rect 197654 70 197854 856
rect 198022 70 198314 856
rect 198482 70 198682 856
rect 198850 70 199142 856
rect 199310 70 199510 856
<< obsm3 >>
rect 2681 987 197603 199681
<< metal4 >>
rect 4208 2128 4528 199696
rect 19568 2128 19888 199696
rect 34928 2128 35248 199696
rect 50288 2128 50608 199696
rect 65648 2128 65968 199696
rect 81008 2128 81328 199696
rect 96368 2128 96688 199696
rect 111728 2128 112048 199696
rect 127088 2128 127408 199696
rect 142448 2128 142768 199696
rect 157808 2128 158128 199696
rect 173168 2128 173488 199696
rect 188528 2128 188848 199696
<< obsm4 >>
rect 34651 2347 34848 199341
rect 35328 2347 50208 199341
rect 50688 2347 65568 199341
rect 66048 2347 80928 199341
rect 81408 2347 96288 199341
rect 96768 2347 111648 199341
rect 112128 2347 127008 199341
rect 127488 2347 142368 199341
rect 142848 2347 157728 199341
rect 158208 2347 173088 199341
rect 173568 2347 183389 199341
<< labels >>
rlabel metal2 s 846 201156 902 201956 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53378 201156 53434 201956 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 58622 201156 58678 201956 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 63866 201156 63922 201956 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 69202 201156 69258 201956 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 74446 201156 74502 201956 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 79690 201156 79746 201956 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 84934 201156 84990 201956 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 90178 201156 90234 201956 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 95422 201156 95478 201956 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 100758 201156 100814 201956 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6090 201156 6146 201956 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 106002 201156 106058 201956 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 111246 201156 111302 201956 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 116490 201156 116546 201956 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 121734 201156 121790 201956 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 126978 201156 127034 201956 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 132222 201156 132278 201956 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 137558 201156 137614 201956 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 142802 201156 142858 201956 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 148046 201156 148102 201956 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 153290 201156 153346 201956 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11334 201156 11390 201956 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 158534 201156 158590 201956 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 163778 201156 163834 201956 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 169114 201156 169170 201956 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 174358 201156 174414 201956 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 179602 201156 179658 201956 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 184846 201156 184902 201956 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 190090 201156 190146 201956 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 195334 201156 195390 201956 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 16578 201156 16634 201956 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 21822 201156 21878 201956 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 27066 201156 27122 201956 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 32310 201156 32366 201956 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37646 201156 37702 201956 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 42890 201156 42946 201956 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 48134 201156 48190 201956 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2594 201156 2650 201956 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 55126 201156 55182 201956 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 60370 201156 60426 201956 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 65614 201156 65670 201956 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 70950 201156 71006 201956 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 76194 201156 76250 201956 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 81438 201156 81494 201956 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 86682 201156 86738 201956 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 91926 201156 91982 201956 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 97170 201156 97226 201956 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 102506 201156 102562 201956 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7838 201156 7894 201956 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 107750 201156 107806 201956 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 112994 201156 113050 201956 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 118238 201156 118294 201956 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 123482 201156 123538 201956 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 128726 201156 128782 201956 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 134062 201156 134118 201956 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 139306 201156 139362 201956 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 144550 201156 144606 201956 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 149794 201156 149850 201956 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 155038 201156 155094 201956 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 13082 201156 13138 201956 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 160282 201156 160338 201956 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 165526 201156 165582 201956 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 170862 201156 170918 201956 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 176106 201156 176162 201956 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 181350 201156 181406 201956 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 186594 201156 186650 201956 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 191838 201156 191894 201956 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 197082 201156 197138 201956 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 18326 201156 18382 201956 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 23570 201156 23626 201956 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 28814 201156 28870 201956 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 34150 201156 34206 201956 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 39394 201156 39450 201956 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 44638 201156 44694 201956 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 49882 201156 49938 201956 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4342 201156 4398 201956 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 56874 201156 56930 201956 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 62118 201156 62174 201956 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 67454 201156 67510 201956 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 72698 201156 72754 201956 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 77942 201156 77998 201956 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 83186 201156 83242 201956 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 88430 201156 88486 201956 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 93674 201156 93730 201956 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 98918 201156 98974 201956 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 104254 201156 104310 201956 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9586 201156 9642 201956 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 109498 201156 109554 201956 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 114742 201156 114798 201956 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 119986 201156 120042 201956 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 125230 201156 125286 201956 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 130474 201156 130530 201956 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 135810 201156 135866 201956 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 141054 201156 141110 201956 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 146298 201156 146354 201956 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 151542 201156 151598 201956 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 156786 201156 156842 201956 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14830 201156 14886 201956 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 162030 201156 162086 201956 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 167366 201156 167422 201956 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 172610 201156 172666 201956 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 177854 201156 177910 201956 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 183098 201156 183154 201956 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 188342 201156 188398 201956 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 193586 201156 193642 201956 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 198830 201156 198886 201956 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 20074 201156 20130 201956 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 25318 201156 25374 201956 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30562 201156 30618 201956 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 35898 201156 35954 201956 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 41142 201156 41198 201956 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46386 201156 46442 201956 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 51630 201156 51686 201956 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 198738 0 198794 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 199566 0 199622 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 188250 0 188306 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 133510 0 133566 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 156602 0 156658 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 199696 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 199696 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 199696 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 199696 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 199696 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 199696 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 199696 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 199812 201956
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 102013146
string GDS_START 1598058
<< end >>

